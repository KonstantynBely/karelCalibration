��  ë�A��*SYST�EM*��V7.7�077 2/6�/2013 A�Q  �����ABSPOS_G�RP_T   � $PARAM  ����ALRM_RE�COV1   �$ALMOEN5B��]ONiI �M_IF1 D� $ENABL�E k LAST�_^  d�U��K}MAX� $LDEBUG@ � 
GPCO�UPLED1 �$[PP_PRO?CES0 � �y1��UREQ1� � $SO{FT; T_ID��TOTAL_EQf� $,NO/�PS_SPI_I�NDE��$DX��SCREEN_�NAME ^�SIGNj�|�&PK_FI� �	$THKYޠPANE7 � 	$DUMMY�12� �3�4��+�ARG_�STR1 � �$TIT�$I��1&�$��$�$5&6&7*&8&9'0''@�%!'�%5'1?'U1I'1S'1]'2h"�GSBN_CFG�1  8 $�CNV_JNT_�* �DATA_C�MNT�!$FL�AGSL*CHE�CK��AT_C�ELLSETUP�  P� HO�ME_IO� }%:3MACROF2�REPRO8�DR�UNCD�i2SM�p5H UTOBAC�KU0 � ��	DEVIC#T�Ih�$DFD��ST�0B 3$�INTERVAL��DISP_UNsIT��0_DO�6�ERR�9FR_F�a�INGRE5S�!Y0Q_�3t4C_WA�4�12HG�X_D�#	 d� $CARD_�EXIST�$�FSSB_TYP�i� CHKBD_[SE�5AGN G�� $SLOT�_NUMZ�APR�EV��G �1_�EDIT1
 �� h1G=H0S<?@f%$EPYO$OPc �0LETE_OKzB{US�P_CRyA�$�4�FAZ0LACIwY1KR�@k ~�1COMMENy@$DGV]QP�� ���AL*OU~�B , $�1HV1AB0~ OLz�UR"2CAM_;�1 x�f$�ATTR��@0A�NN�@�IMG_�HEIGHyAcWoIDTH�VTC�YU�0F_ASP�ECyA$M@E�XP;$� Mf��CFcD X '$GR� � S!1U`=BfPNFLIC`~d
UIREs3��A�OMqWITCH�}cX`N.0S_d�SG�0 � 
$WARNM'@f��@�� LI? �aNST�� CORN��1F�LTR�eTRAT�@0T�`  $ACC�1"p '|��'rORIkP�C�kR�Tq0_SF� �!C�HGI1 �[ Tz`u3IPpT�YVD�@*2 �P`�`� 1zB*HD�SQJ* ��q2�v3�vU4�v5�v6�v7�v�8�v9�E �CO�$ <� so�o�h��s1�PO_MOR~. t 0�Ev�NG�8`TBA� 5c���A�����]@����ϋaP�0Ѕ*��h�`
P�@�2� �,p�J,p_Rrrqo@+�1J/r/�J�JVq@��Cj��m�g��ustP�_}0OF� 2  @� RO_���Wa�IT8C��NOM_�0�1ەq34 ��cD� �;����hP���mEXpG�0� �F�p%r
$TF�x�JF�D3ԐTO��3&@U=0�� e�H�24�T1��	E�� �e��f���f��0CPDBG�;a� k@$�PPqU�3�f):�L�A�AX 1�dUN�v$AI�3BUFuF8����! |�`��`PI��P�r�Mq�M~�䠁�F>r�SIMQS���G��QE������MC�{� �$}1JB8�`S�}1DEC���������x� ě0CHNS_EMP�rG$Gg�=Ǎ@_��<q3
p1_FP󔞡TCh�@`�b��q0�c}�y�G�� V�AԂ�!�!���JR!0ԂSE�GFRA.pv 7aR>�T_LIN�C��PVF������Y���Q��)B|����( '�� �f�e�S���Q��.0��p�B��A����SIZC�ћ�z�T��g���|���QRSINF3� �p����?�������؄����Lot��G�*�C3RC�eFCCC�`+� ��T�h��mh�SbA�� h�*�f��:�D�d�c2��C��PTA����0w@�撀��EV���jUF��_��F��N&��G�� X����r��1i��! ���,��hRGNP��0qF����R}�D���2}�LEWN��Hc6���C��K�۲RcDx :�L��ou2���A6uN`Co�$LGp��B�1aP��s@�dWa!A?@���~0R���dME%`��d�_3RAs3dAZC�4��z�OkqFC�RH`�X`F�`��}��,�ADI;� 6b� ����`�p�`5cn�S0�@1�7a�AMP���PIY8CU�MwpU��:iQU� $�P���C�CG1������D�BPXWO����p$SK��2��wDBT TRL�1	 ��Q0Ti� �P��DJ�4LAY_C�AL�1R !'P1L	3&@�0ED�Q5'�Q5'̡����1�!�W�PR� �
�1 0�1" l�PA$�q$��/ �L�)#�/�#�mp�0$�/�$C�!%��/�$ENEqr�1&�/�#d REp�"_'H �O)@o"$LF3#$�#�xB� W;���FO[ _D0m�RO(@���u���j���3RIGGER�6PA%S��ETURN�2RcM[R_��TU�`?�u0EWM����G1N�P��zBLA��E^��$$P#�CPD� ��&@�Qk�C5D�mpD�A#�p4\1i���FGO_AWAYF�2MO��fQg�wCS_(<�QIS ����c�C���A����B�t�C�n��A"�FW���DNTV@��BVkQ���� �S˳W�sU�J&�U�<� ��SAFE�ZV�_SV6bEXCL�Ul�����ONL�A��SY��Q�tOT<Ba��HI_V/M�PPLY_�a��VRFY_#�q�Bd�_ )0���9_+�Ip !��A;SG3� *�b݀ �0 AM���a*����0ⰀVi.b%fANNcUN� rLdIDp�	U�2~S@�`mija�rj�f�RpOGI:�"+��$FOb��׀OT@w1 ?$DUMMY���d�[!�d١�& �E,o ` 8�HEx�s��b�SB$�SU7FFI�@ ���@�a5�g6�a.��MSW�E- 8���KEYI����T�MZ1^ӌq�1�vIN������. �D��HOST? !�r���t[ �t٠�tYp�pEM>���$���SBL��UL��/� �|3����T�50�!0 � $<9��ESAMP�ԕ F��������I�0�>�$SUBe�Q��� �C�:��G�SAV��r���G�C� ˇ,�PnfP$80E���YN_B�1 0&��DIad�@O���v}$]�R_I��� �ENC2_	ST � 2
ԇ J���L�q~S�`;����!!3�M�I��1:�p�4  L�3�M���0�0K�4'a��A�VER�q��}�M�D3SP�v��PC�U����\ì�VALMUŗHE� ��M�sIP@���OPP7  �THS ���6��S�F�F􁳠d0L�0�T��SC�Q�dm:�ETo�5zrFULL_DUY��da�0��O�w�h�O�T���0NOAUkTO�!6�p$�H\���cl�
�C!�e�C���"���L�� 7H *�L���n�b���$�0P�˴��ֲ�� [!���a��Yq��dq��U7��8��9��0�����1��1��1��1�Ⱥ1պ1�1�1J��2
�2����2��U2��2Ⱥ2պ2�U2�2��3
�3���3����3��3Ⱥ3�պ3�3�3��4�
�[���SE�"8� <��~��`�;I`�����/��QFE�0��0� 9 ,��Q?g z@^ ?��А��ER@#�� ��@��� :�`$�TP�$VARqI�<��UP2�P3; �pq�TD��S�|�1`3���qr�B;AC�< T�pr���)��bP��@o�IFI)�@���U���P��F�0��� =t ;'�Ԡ��P'�ST(&�� HR&�Pr0E����	%�C��	���_Cr�N�r��B���p�h�FORCE�UP%bn�FLUS
�`HN �E�h�R/D_CMK@E(����IN_��&vPg�REMM�F~Q���M �� 3
K	N0�EFF��N@sIN�A��OVMl	�OVAl	TROV̙��DT��mDTMX���m{@�
���? �*[ ��CL���_:p']@$�-	_�
�;_T��X
�J�@AQD� ��}���}!V1� RQ~��LIMIT_�ad椀�M��CLmd�}�RIV	�a��E�AR��IO*PC�C�����B�Bg�CM�@��R �GC3LF�G!DYM(/l�aR#5TWDG���| s%�+�FsSS& �s> P�a(�!r1��wP_�!�(J�!1��E�3�!3�+=5�&�GRA����?w��kPW��OyNT��EBUG)S�&2*�P{@a�_E �@�P�Q@�T�ERMB5AK5���ORIG0BK5 ?�
�SM_�Pr��G0C{6�PTA�9D�K53��UPB�Eg� -zAa�@.P|Y3.@A$SEG�:vf ELEUUSE�@NFI,��2�1xޠp4�4B$UF6P�$�FQ4@�wAG0TQ�&�HSwNST PATm�<piBPTHJ�AߠE�p��2�P؀	E)��؁��1R�@�InaS�HFT_��1oA�H_�SHOR ܣ�6 ��0$�7�@Dq�'�O#VR#�na�@I�@��U�b �QAYLO=�z��I'"�oAj�!�j�ERV��:Qh� �J��OG @�B0����U�>���R!P"�AScYM.�"��1WJG�уES�A�YvR�U�T @���E)�ᥳEaP!�WP!�WOR @�MB��GRSMT�F�GR��3la�PA.@��`�q�uG� � ����T�OC�1�`P�@ �$OP��ဝpՓá� ��O��RE�`RC�AO�pтpBe�`RmE u�h�A���e$PWR�IM�ekRR_�c4��q.B H2H���p�_ADDR��H_LENGqByqnq�q��R��S�I H��S���q0Ӧu>Ӵu���u��SE�'�LryS��J $J�<�`��_OFF��r�PRM� ��HTTP_�H��K (^pOBJ�?"ip��$��LE�`C!�ȠL � ��׬�AB_~T�S�s�S{`��*�LV�N�KR��eHIT���BG��LO�q t�fN�͂���`���`3SS{ ��HW��A��M�p`INC�PU�"VISIO �����+��t,��t,�~�� �IOLN���N̠�C��$�SLQb��PUTM_�$�`{�P x�V���F_AS�"O��$L��I���D�A��U�0�@Af��`q�<PHY���Ó̞1��UO��#P `������ڔ� �2�pP���`(�L��XY�B��!UJ�Q�vz�NEWJOG-GN��DISx�[�K-�Lf�#R 
�WAV��ǢCTR�CǢFL�AG�"[�LG�dS� ���Y�3LG_SIZo�����X����FD)�I� 4�E�*��D0���c $���𖶦���K���xD0��� SCH_���߅p�2��N��F�T
���E�"~�����"��U
�
�{`L�	�7DAU/�EA�-��dE�;�GH�b��BOO��Uh Aɒ��IT��y�[0�ŖREC��SCRX��ʑDIēS.@��RGO���˒�����d�´���SU���Wp�Ĳ�Ľ�JGM$��MNCH,�FN�KEY%�KM�PR�GK�UFY�PY�F�WDY�HL��STPY�VY�@Y؀�Y؋RS��H1`uۺ�C�T���R��� �$�U 	�m���
R�ݠғ`�G=��@POd�ڻ�z��M�FOCUd��RGEX��TUIK�I{�����	��� ���I�M��@A�S���`���@������AN�A���2�VAIL�l�CL!�UDCS�_HI+4`�s_�O�e�
!h�S���|�S����IGN4��F��J��T�be�_BUTj � V !PT�$*��rv�Ϥ�(���a�!W !Pi�P'���0�1?2?�3?��_� X � i�=a�5����&��ID� tbP5R�baOh ��\A�ST	��RF�Y� �@�  /W$E�C�y�����_�� Y L�؟0��@�� �`qFtǀ�FwҬ�?_ Z �p�����b���>0C��[{ �p CLDP	�>�UTRQLI{��T8����FLG��� 1�O�D�����LqD���ORG�� ����hW>(�siT�r� 4\ �#0��Ք��Sy`T�70�y ' �$�!�#RCLMC�$B/T/�)Q��!r=1I�p_d] d��RQ73$DSTB�p�   6��-8�AX�R /8I<E�XCES�b�12Mp�1^��2�Tt��2��0_�p"6_�A:&��;G?Y80K�d` \�GRO�U��t$MB �L�I9�CREQUI�RDB�aLO#KDESBUr�u1LYM���agbʑ`@�C�"Fu1ND��`c`b��̨�CDC���IN'��C��Z`���H��N��a#�� �EP�ST�� c\rLOC�RITp��PAp�1u1OD�AQ��d X�O	N�cF�R�fV�	�X��b�U���w ��FX0IGG�� e �y X�a��hX�XR�Q%���Y	��X	��V�0ғD'ATA$`E�a���a�N��f t �$MDEaI:�) Sf��^d�![gH5P�@�]ez��a_cANSW��a^d�a��^eD�)pARz�� Xpg �0�CU4�V�`�=UR;R2{�h D2�`A���A�! d$C'ALI&0��GS�w�2K�RINb�t<N�NTEg�(i�b`Cu��=RBqg�_N�q�jPukr���$ht�2knuyDIV�&DHi0tjp+�l $Vp�C�$M�$Z 0R<!T 0R���b�e�mH �$BE�LT˪ZACCE�L���;�"�IR!CO�݁m��T���O$PSi0�Lt0ڰW��Cp8��T�9�PATH���.�"��3]��Pl1_<�r���Ł�"S Cr��_{MG��$DD�<9���$FW�`7``���.���DE��PPABNe�ROTSPEEՂ@L� JN�@��(0�t0?$USE_p�P&�ܦSY>��p�!- �QYN0A�����OFFua��MOUf߁NGJ�܀OL~�ٔINC�d2Q���-2��� -2ENCS�pa2U��+4R�IN�I]�B����"n��VE��s^�23_�UPօp�LOWL���[�` '���D�>�2@Ep]'��2C�[pW�MOS���4M�O��0�'PERC7H  ��OV���� 蓼������$�8S@+�� 2@������V�0^�O�L�P��7O��U�UP"�������T�RK��AYLOA�J��1��]�͵³83P� �RTI�1	�� MO�O�-2�28 �`4�wٳ��?��pDUM2��S_�BCKLSH_C ]�P�ϐΦ����bn��"�y�Ñ���CLA�L V��!��� ��C�HK �SՐRT�Y����C�
*!6a_��ä_UM����C����SCL�W�LMT_J1_L< "0-օa:�E4�U��G�D�J�P�J�SPC`d�ȑZ���3�PC �B3�H_A@���C� �cXT���CN_"rN���.�S��%�V���:����]�d9���C' �SH� r�*�*!9�9� p��0^���9���PA���_P��_�"�Ŷ`�!ճ����JG�����~�OG��,�TO7RQU��ON��޹�*�B٢-�*�L�_Wž�_�sj��sj��s�j�Ir�I��I�sF�KP]�J�!��c!�VEC�0'42��1��p{0��82��JRK���+� DBL_S�M���"M�@_DL�q�"GRVq�j�sj�sKH_��I����
COS��LN- �����p�	�p@�	�����FZ� �٦KMY�D�T�H�eTHET0��NK23�s��s�� CB�CB�sC &1n2�����s���SB�s��GTS�1W�C.�2Q������$�'3$DU ���8A!r�2P&�r1Qb8V$NE�4��PI� ���"%�v$�p�A��%�'���LPH�5�"h��"S��3�33�"P+3:2�pV�(V�(T�p�,V�*V;V;UV";V0;V>;VL9H�(�&�2�-n�H;UH;H";H0;H>;UHL9O�,O�(O}I��.O�*O;O;O�";O0;O>;O2F��"�Y�T�'SP�BALANCE_lT@SLE�H_�SPHq�hR�hR3PFULClX�R{WؓR3Uz1i
�UT�O_����T1T2�Y�2N���`��T�q���Ps d���T��O�p!�L�INSsEG���REVf���Q�DIF��zy1�j_g�r1k]�OB0Ua��t$yMI`���~SLCHWAR>���AB��u$MECH�Tˑ�a��AX˱Py��f�'�r�Pl 
�bI��:�7ROB�CRW�-u��ҏ+�MSK�_KP�tn P 
�P_��R��r_tn���18�c�a�_p`�y��_p�aIN:a�M?TCOM_C���po  ݀g`4�?$NORES��ry��`�rp 8U�GRJ��eSD?�A�Bג$XYZ_�DA�!F�r�DEBaU:a�q���pq _P�$��COD�� �1����`��$BUFINDXa�w  !�MORRs/r $�qU&��ƀu��ӑy�W�!��bG�i�s � $SIMUL��8��>�<��F�OBJEjP���ADJUSψA'Y_I��8�D����s�Ԑ_FIב=s�TZ��c����`@b�"�(�b`p0G�D���FRIW�d�Tg�R�O%�A�Eb�GqO�PWO> Vpt0>>�SYSBU0[�$SOP��I�����yU��b`PRUN�rڕPArpDٖ�b��.1�_OUTΑ�a��t$�IMAGҊ�\pv PDaIM���1�IN[ �0�RGOVRDY�˒����P�/�a�� L_`�PB�}����RB��s���MkᜪEDTb��` �N�@M��2~�^�\�SLjPVp�u x $OV�SLfSDI��DEX���q�����o��Vb��N�A�� '��,�'�D�M~]��ӣ_SETK�Vpv� @U�^��ep�RI��j�
q�_�}����^�dà*� �w H\q�`��AT�US<�$TRCpx T�X�ѳBTMڷ*ıI��P�4}Ѱ�\��Vpx D\pE���β�0Ehbϱ�����ϱEXEհ����)�=��f�ym�]p԰3UP�L�$�`6�XNN����������� �PG�uzWUBñ�e��ñ���JMPWAI[�PL���LO7о�FA`���$RCVFA�IL_Cwq����R 9��p�c��(�}�"�-��AR_PL��DB�TB��,⾐BWD� ��pUM*�"�IGp�7��Qc�TNLW�D"�}�Ry�iӻ�E�����^���DEFS}P` { L\p��`��_��Ճ��UN!I����Ѐ�RD��R�b _LA`PͱY�P�pUq|-�#��q�O���XPc�N�PKET��
��Pq�Uq}� h�ARSIZAE5p��=��u�S̀�OR��FORMAT�Pg�COנq�<b�EM�d����UXx��,����PLIb�~Uq~  $�p�P_SWI�`���^�/ G�b�AL_ So���A�rB���C�rD��$E6L���C_lі� � � ����r��J30 �r��TWIA4Z�5Z�6�rMOM��f��s��4��pB��ADf���s����PU�NR ����s�������Rt��� A$PI �&E�kqE�p-~- �-�WC�0$���&�9q�gE��eS/PEEDL@G�� ���Ծ����)�9�����)��	)���SA�MWPx�0�1��MOVD�H$_S`Y%nHk%_��1�t�2�t@����c�v��8�H�PxIN����������(�+(+G�AMM<Vu!�$GGETE�U�ٓD5�z��
�PLIBRv����I�$HIu�_�L�ݰpB�&E�(A�.� �&LW�-�&�, �)	6�&1��f�`j���� $PDCK���ٓ_�����E���b7��a4���a9�� $I��R�`D�c�b~�Ե`LE�qkq���8�1��0�Gq��`Vp��P/aUR_SC�R��A�r��S_SAVE_D��8Ex�NO5�C��y�6�8@ {$E�.{I��G	{I�@ �J�KP�q��H� � ��x"Mao���s ����d��6W2U�C�qy�����M� �k�F��aE��3�W<�@[�jQWg@5r�U��R�R��Sc2jQML"��[CL�W��M)A�Tr� � $P9Y����$W`�fNG�O�`�b� b�b#�HЈ��a� (���c��X�O����Z�e��ހRt� p䠰p�3+zO�O�OаO�O�a5�_�r� |�E�8@��>vs�>v@��8@_�kwVvy�Eހ�u% ��"rB��\�P�"tP���P�M&�QU5 �{ 8*�QCOU�1QTH#pHOL�<�QHYS��ES�e�qUE�p.BZ�O.��  q�P���%杲UNְ�Q r��OE��p� P2��3��AÔ�ROG(�����Q2(�O}�2�x�����INFO�q�� #�e����R�v��OI��� (�0SLEQ�с�рHi�C�{�D��L��`�� OK0r��!E�� NU!��AUT<TA�COPYqu�(?��`@ML�NI�M��X�Cᐛ� Y�RGWADJ�q�i�X�Q���$ഖ�`��W��P���0�������[EX8�YC0b�ђ�Obp�q���$�_NA9!��������`��� � 9Q���POR�A�\B�SRV0�)a�6Y�DI��T_��{��������������5*��6��7��8y����S8BL��m�MC_)F�p��PL9A8An�ȰR��9��Ѽ���$iB����d� ,ƨ0FL-`L�C@YN��[�M��C?��P�WRc��L��!�D�ELA��8Y5�A�D�a���QSK;IP� �Q�4�-OR`NT�� ��P_4��ַ@lbYp �������� ��Ƞ��ՠ������z��9�1�J2R� nL�� 4*�EXs TQ%����(Q�����p�����p���RDCNf� �`��X9�R�p�����r��A$�RGEAR_� I9OT�2FLG��vi̥�M%PC��B�UM�_����J2TH2yN'�� 1������G8 T00 �$����MlѺ`I�8� REFr1�q�� l�h��ENAB{�(cTPE�0�1� ���i�m���^QB#��@:��"������2�������������&�3�Қ7�I�[�m����&�4�қ������P�����&�5�Ҝ1�@C�U�g�y���&�6�������������&�7�Ҟ+=Oas�&�8�ҟ������&�SMSKJ�q�|��a��E?A���REMOTEF����a@��L(Q�IOQ5�Ic:(P	��POW�0L�� �pZ����#p�%�L��U�"$DS?B_SIGN�1)Q�%���Cl�(P��S�232��b�iDEVICEUS�|,R'RPARIT���D!OPBIT`Q�Y�OWCONTR`;�(Q��O'RCU� �MDSUXTASK�T3N�p[0�$TATU`PV"�0L�����p_,PC9��$FREEFRO�MSp��%�GET\�0�UPD(�A�2�V"P� J���� !)$USA�^���6���ERI1O�P@bpRY�5:"�_>@ �P}1�!�6WRKI[D���6��~aFRIENDmQ�P$UFw���0oTOOLFMY�t�$LENGTHw_VTl�FIR�`�-C�RSEN ;IUF�INR]��RGyI�1ӐAITI��b4GXӱCI�FG2�7�G1��Ѐ3�B�GP1R� A�O_~ +0!�1REЀ�E3ⅆe�TC���Q�AV ��G8��"J��� u1~! ��J�8�%��%�m��5�0G4�XS _0)�L|�T�3�H6��8���%r4E3G�U�W�P�W�R�TD ����T��а��Q�T�m�$V 2�����1���91�8�02*�;2/k3�;3�:i va�9=i�aa�^S��jR$V��SBV�EVP'�V�BK�����& c�p��F�"{�@�2�q�PS�E��$p.rRC��o$AŠ�FwPR��Gv]U�cS�'�� 7�6A6I��# 0�@qV`��p�d�`���E0�@��=�
zB5S!� ��a�Rg����R�6�N� AX�!$�A�0Lx(A���rTHIC�1�Y���h�t1TFE�I��q�uIF_CH��3�qI�G�a�pG�1bxf���m���S@n��_JF��PR��ֱ�S��Ԁ�d� �$SР�Z�G�ROU�̃TOT��t̃DSP�JO1G���#��_P��"�O�����j��&KE�P(�IR����@ML�R@�AP�Qn�E^�8`�!�[�SYS6��"v[�PGu�BRK�B( �.��pIq�p��0M���΂�`AD�!̃�9�BSOC׆�N�ӕDUMMY14�p@SV�PDE_�OP�#SFSPD�_OVR=���C����OR�CN�m0�F.����OV���SFR��pU���F�n��!#��C��A�"LcCH����РOV�s0��W�@M��ĥ:�#RO�#ߑ�_�p��� @@�u@VER��ps0OFSu@CV? �2WD6���2�ߑXj2Y���TR�!����E_FDOY�MOB_CM�D�BBL�b>�f��attV@"Q�240/p��N�Gg�z�AMx�Z�0���¿_M~��"7����O8$CA�7�D����HBK81���IO�5���QPPA�=�"�M�5�͵����DVC_DB xC~� �3"�Т�!��1��糖�3����pН�*��U�3��CAB��2VӆPѣhIP��c�O��UX�?SUBCPU`�	�S�P P���90^SQ��c��."��$HW�_C�Т��S��cA��A�pl$UNIT���l��ATTRIx"���	�CYCL���NECA��J�FLTR_2_FI_�0G(��9&�1LP�?��>�_SCT�CF_ƣ�F_��6��FS88!����CHA�1�pwᇲ�"v�RSD�`4"���a��_T���PRO��>�� EM�y_ܠ��8d��ac d��a��DIb0~!�RAILAC��9RM��LOÐ C딂�Q*q��3q���P�R��SQ�pU�C�r�s 	�FUNC��@rRIN'PѸ0���u��!RA��B �����F�Ğ�WAR~���BLQ����aA��������DA��0��	����LD)0���Q1�q��*q1TaI2rQǁ�p$xPgRIA1�"AFB�P�!|ߠ�<`�R����MOI��A�D�F_&@��51��LM���FA�@HRDY.�4ORG6 H���A��0 �MULSE�&@"�Q��a �hG�	�����$d�$�1$1 ����0���� x�m�EG�̃�`A1Rހ��09�2o���z�AXE�RO%B�W�A��_�œCSY������S�'WRI�@s1�ЇSTR�� ��(�E�� 	%1��A�B( �/&�a�ӰO�T0^�	$ߠA�RY�sf"���S@	��FI��*�$LGINK���!�aI_%#�%{q�"�XYZ82�*�q�#O�FF���"�"�(j B�j�4С��n�3FI��%7�q���j���_J���%���#�QOP_>$H+5��3�PTB\1�2CL��i�DU�&62�TURN��2r�5t!0}��p��|7FL�`�� �m�0�%+*7�	�� 1�. K�M�&82�Q�2rQ�#�ORQ��G��-(� +p��z�� 3q�E"�T�GOV�@-A��M *�y�4�E:�E@�FW�J��G���D��o� *� ��A7�P��y� �E�A�GZU:ZU�CG�SER���	6�E���B�TAFQ��)4��`��r'�AXУ a2.q�c�W�c�W�c �W�p�Z�0�Z�0�Z%@ �ZK@�Z��Z
!�V�  �Y� 
i� i� *i�  :i� Ji� Zi� ji� xzi�a�iDEBU{�$v�u��;q��"F7O�n�AB��6�r�CV�z� 
fr ����ukњw�!�w�! �w�1�w�1�w%A�wKA��w��\0��"3LAB"2|EwЄ�҂��3 � EER�VEN� � �$q�_NAǁ!_�PO����` f��M�_MRA��� �d  T���EcRR����~ TYi���RI�V"0�S��TOQ�T)PL��T��Ѕ
L�G�CJ � p�PTl X���_V1�b�Q���#��2�2+�����/@�8�p��5�$W��V�j��VN�[�$�@@�� �S���Q�	E�HELL_CFG�N� 5%�Bo_BAS��SRvp\0�K� �S��TJϐ1a�%Α2�U3�4�5�6�e7�8�RO࠘��� � NL:�3AqBn��АACKwv ��)�o�u0iႩ7_PU2�COq��OU��P��ӕ������TP�_KcAR�0��REm��� P��z QUE�٩��@���CST?OPI_ALzs���� �TĠ�� SE�M[�w�k�Mw�y�T�Y��SO`��DI����Є�=�װ_T}MK�MANRQζ� E��$KEYSWITCH���Ѱ��HE��BE�AT��R�EpLE(����&�U��Fd���|��SO_HOM� �O��REF�@PR�i��R� ��C@�O0�p ECO���� _IOCM�4M�k��^����'�O� �D�!ۧH�U��;�M�7��@�3FORC�ߣ�� ��OM>q � @Etx*k�U#Po1B�O��o3B�4x��N�PX_AS��� �0ݐADD��(��$SIZߡ$VsAR�TIPr�)q�G�A(ҷ��
� ˨r�t�n�SV�XyC����FRIF�R�S%�7�x���NFpѲEАO� x�PSIڂTEC*�%C�SGL=�T�"�0&��V�D��>�STM�T
�o�P\�BW<�@?�SHOWw��P��SV� K��; ���A00�0�Q ��K���O���_���iЪ��5��6��7��8
��9��A����6� �����20��F��
  ����U ����� ���@�0�� �J@��:�1G�U1T�1a�1n�1{�U1��2��2��2��U2��2��2�2�U2 �2-�2:�2G�U2T�2a�2n�2{�U2��3��3��3��U3��3��3�3�U3 �3-�3:�3G�U3T�3a�3n�3{�U3��454��4��U4��4��4�4�U4 �4-�4:�4G�U4T�4a�4n�4{�U4��555��5��U5��5��5�5�U5 �5-�5:�5G�U5T�5a�5n�5{�U5��656��6��U6��6��6�6�U6 �6-�6:�6G�U6T�6a�6n�6{�U6��757��7��U7��7��7�7�U7 �7-�7:�7G�U7T�7a�7n�7{��7���VP$�UP}D��  �Px���x�YSLO��� � ��հ�����QTAS�sTƠ���ALU}U����C�U��WFdQID_YLѳ�UHI�ZI�?$FILE_Σ�Tf�$u�_VSA��� h��+`E_B�LCK(�8bg�AhD_CPUQi��Qi����Sod_R1�ɢR ;��
PW,�d�[ �aLA�S��8�c�a�dRUN5��a �d�a�d��5��a�d�a��d �T�pACC����X -$&qLEN~�3t��&p䫠��Iѱ
�LOWo_AXI(�F1&q
�T2mwM��ɢ���I����Q�yTOR.�&p�{DW��s�LACE���&p�����_MAuйv�u�w�qTCV�|��wTڱ�;�1�<ѷt��H_��s��J����M��"��J����u���u2q2��������s6�pJKцVK~��4���3ՃJ0����JJ�JJ��AAAL�����4�5Xr;�N1B�N��	��tL�p_k��nѼ"p��� `5`GGROU�PY�ӲB$ПNFLIC�ө�R�EQUIREv�E�BUV�"q���кp2����#pɖ!qxг��� \��APPR�ՐC���p
!�EN��CLOz�,�S_!M ���A��u
!q��o� 䣠MC�r8;�Xr|�_MGц��C��,`��N��p��B;RK��NOL����:��Rϰ_LI��է$����JޠѤP��p ��p���p;��pD��pQ6�K��8��/��>���� ҒMr�:ql�Gqz�PATHv�������Rx��������pCNR�CA���է���IN%rU�C�pwQ�Cd�UMB�Yop�����QE:p��Gp�����PAYwLOAͧJ2LHPOR_ANqQ�L�`�[�W�K�g���R_F�2LSHRё�L�O\�䱕����ACRL_�����޷�C�XrH�P"�$H����FLEX�� qJ%u� : 2Dv�p4�K�GYq�pPbt|F1Kљխ׀��������E ����/�A�S�e� w�����y���ф���� ������J�ÊT���X����υ ��څ�� [����
�� �)��@;�D�V�h�z�Y�J��� � ��������QIPAT��ё��EML4� �ؘJ����ߐJE��CTR,ޱ��TN��F�ɗHAND_VBp�qѹP`�� $&��F2��K��ШRSW�q?QTBj���O $$M��}�R���E��Uw�H��sA@�PH����Q���A���P��A��Aɫ���Tj`��D��DɫP��G�`1)ST��9!��9!N̨DY�`��� |�Y�鰋�KыǦ�@J�ч�s�U�ХP� �&�/�8�A�J�S�=��� ; �t�.Rx66N�/QASYM����Ґ����Խ��ٿ_SH�����筀�4��+�=�O�J�V��h�'CI����_�VI�dHN�u@V_UNI�ÉD���J҅�B�%�B�̦D�� �D�F�̓�������τ*Uc���X��H̴`��XQENL� v�DIɠS�OwTqY�YP��� ��
�I�1A��äQ�`�Bc�S`�  p�a.a�o � ME����R'R�1TkPP�T�0) ���Qz�~� ��0�Xa	iT@�� $DUMM�Y1��$PS_6��RF��  ��Pfm�aLA��YP��jb�S$GLB_T>mU�e�PpQ p���Q� X	�ɗ`��ST��ߐSBR���M21_V��8�$SV_ER��O�Ð�c�cCL�`�bA�5�O�RTPT O�P �� D �`OB���LO˰&uq�9c�`r�0�SYS�qADR�TP�PT�CHb � ,x&����W_NA��c�tz�9SR��?�l =�� M�u`�ys�u~�s ��s�������� ���0�)�T�"�5� ~���B����s�?�?�?|DY�XSCRE)�jp�ȐST[�Fs}�P!��t)�r _� Aq� T 	��`ob��a`�l��Ҩ���g�c�O� I�S�c��T!Y�UE�T� �ñjp^`ySq�RSM_iq�mUUNEXCEPlV֑XPS_�a�����޳����޳R�CO�U�ҒS� 1�d�UE�tҘR�b9��PROGM� FLރ$CU�`POX?Q�д�I_�PH��� � 8џ�_�HEP�����PRY ?��`Ab_Ѹ?dGb��OUS�� �� @�`v$/BUTT�RV`��COLUM��U3��SERVx��PASNE� q��P@'GEU�<�F���q?)$HELPB�l2/ETER��)_�� m�Am���l���l�0`l�0l�0Q�INf���S@N0�� ǧ1�����ޠ �v)�LNkr� ��`rT�_B���$H�b TEX�*��ja^>�RELV��DIP�>�P�"�M�M3�?�,i�0ðN�jae����USRVIEWNq� <�`�PU�P�NFI� ��F�OCUP��PRI�8 m@`(Q��TR�IPzqm�UNP�T� f0��mU�WARNlU��SRWTOL�u���3�O�3ORN3�R�AU�6�TK�vw��VI͑�U� {$V�PATH���V�CACH�LO9G�נ�LIM�B����xv��HOSTN�r!�R��R<��OBOT�s��IM
�� gdSX`} 2�����a���a��VCPU?_AVAILeb��+EX��!W1N��=��>f1?e1?e1 �n�S��; $BACKLAS��u�n�\��p�  fPC��3�@$TOOLz�t$n�_JMPd�� ݽ��U$S�S�C6��SHIF ��S�P`V��t�ĐG�R+�P�OSU�R�W�PRADI��P�_cb���|�a�Qzr|�LU�A�$OUTPUT_3BMc�J�IM���2p��=@zr��TIL��'SCOL��C���� ҭ�Һ����������o�od5�?�҂Ȧ2Ƣ�p�0�T���vyDJU2��� _�WAITU���´n���%��NE>u��YBO� ��� $UPvtfaS�B�	TPE/�NEC��� �ؐ�`0�R6�(�Q��� ش�SBL�TM[��q���9p���.p�OP��MASf�_DO*�rdATZpD�J����Zp�DELAYng�JOذ��q �3����v0��vx��,d9pY_���	�7"�\��цrP? ��O�ZABC�u� ��c"�ӛ�N� ��$$C��������!X`X` =� VIRT���/΢ ABSf�u�1 ��%� ?< �!�/ �/??0?B?T?f?x? �?�?�?�?�?�?�?O O,O>OPObOtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo Zolo~o�o�o�o�o�o��o�o{� ��AXL�MT�s��#  �tIN&8qtGPREO��+vup�XuLARMRECOV �)Xrzu�jF �%�!d�� ����7�I�[�m��~�,� �/��uN�G5� �+	 �A   ڏ�� PoPLIC5�?�%�upՁHa�ndlingTo�ol -� 
V�7.70P/36�뀬�
]�_SW�2�D�F0j�W� �43Y�J�9�K�7gDA7?����
&��X�e	-�Non%e��J����� �T7�	���E_�Viu�6s��UTOz"�,tTy.�?HGAPON� %���!.�U��D 1�y� t�x�����xy.�K�Q 1�{S  Hp�������	���uq��"=�" �!���Hեw��HTTHKY��"ٯ� ���u�����󿽿Ͽ �����)�;�M�_� qσϕ��Ϲ������� ��%�7�I�[�m�� ���ߵ���������� !�3�E�W�i�{���� ������������/� A�S�e�w��������� ������+=O as������ �'9K]o �������� /#/5/G/Y/k/}/�/ �/�/�/�/�/�/?? 1?C?U?g?y?�?�?�? �?�?�?�?	OO-O?O QOcOuO�O�O�O�O�O�O���TOĀ���DO_CLEAN�D���{SNM  ɋ���_�_�_�_o���_DSPDRY�R�_��HI!��]@ �_}o�o�o�o�o�o�o��o1CU��MAX �bTQNQS�sq�XbTB�o�B���PL�UGGb�cWo��P�RC4`B�P]k�lo^�rO�r=o��SEGF;�K�+�6� �_�_}�������ŏ�0�LAPZom�/�� +�=�O�a�s�������ໟ͟ߟ�6�TOT�AL�v�y6�USE+NUZ�g� HXL��NR��RG_STR�ING 13�
_�M,�S��
��_ITEM1��  n󝬯�� Я�����*�<�N� `�r���������̿޿���I/O �SIGNAL���Tryout �Mode��In�pB�Simula�ted��Out�T�OVERR~W` = 100���In cycl�Hŕ�Prog OAbor^Õ�>ĿStatus��	�Heartbea�t��MH Fa�ul����Aler �����'�9�K�]�po߁ߓߥ� ^S ��^Q��������,� >�P�b�t����� ��������(�:���WOR9���r���L� ������������ *<N`r���p����PO�� �����9K]o �������� /#/5/G/Y/k/}/�/DEV� -�/ �/�/??)?;?M?_? q?�?�?�?�?�?�?�?�OO%O7OPALT��^A��8O�O�O�O �O�O�O�O__(_:_ L_^_p_�_�_�_�_�_LOGRIxp��avO �_*o<oNo`oro�o�o �o�o�o�o�o&@8J\n�_*�R�� �qo������ (�:�L�^�p����������ʏ܏� ���PREGbNK��$�r� ��������̟ޟ�� �&�8�J�\�n������������$ARG�_r�D ?	�������  	$�W	[�]����.��SBN_CONFIG ���L�K�F�CII�_SAVE  ��k�b��TCE�LLSETUP ���%  OM�E_IO��%MOV_H��¿ȿ�REP�|��UT�OBACK���V�FRA:\8� �8����'`��8�c�,�I�NIa@8�^�~,�MESSAGz��������ODE_!D��}�C���O� ���,�PAUS!�~�� ((O�� J�\�F�|�jߠߎ��� ����������B�0��f�t�%�*TSK � 5ݒϕ�/�UP3DT����d�����XSCRDCFG� 1��� 	�������&�8�J� \�n���\�n������ ����"��F��j |����/e�>2�GROUN��߾�UP_NAܰ���	2��_ED���1
��
 �%�-BCKEDT�-��}��p���g3�p8�/�,/�8���g2���E/��/��/~/��ED3n/&/�/�J/\.�/"?�/�/ED4?�/?�/\.[?�?5?G?ED5�?n?#O��?\.�?jO�?�?ED6ZOO�O6O\.�O_}O�OED7�O�Ok_��O\.G_�_!_3_ED!8�_�o�]-�_8Vo�_�_ED9Fo�_�o"o]-�o�oio{oCRoY_Vh�]1��{� LNO_�DELGE_�UNUSE	L�AL_OUT �V��WD_A�BOR���~�5�I�TR_RTN�ǀ�H�NONS)Ю������CAM_PA?RAM 1�����
 8
SON�Y XC-56 �23456789�0Y �f�@����?�W�( CА��8�h�х�ڎ��HR5ǃ��	���R570�B�Affފ������ڟ �ǟ�"���F�X�3��|���i���į!�CE�_RIA_I��j����F��;��Я ���GP �1�� �s�����V�C󠸾i����CO�C ��Y(��ǀC8��@���H��CCX����C�h��p��x����W C�����Ⱥ���+�=�G��ށ��H}E/pONFIG=��f�G_PRI 1�B�$r�����������(�~�CH�KPAUS�� 1���� ,wuj�|� �ߠ߲���������� �0�B�T�f�x���4��D�O���T���_MORGRP7 2?� �\�� 	 �,��P�@>�t�b���5�����$e�.�?a�a�����QK���d�P�V>��a�-`�/A�

s��� ����b&�i��ܦ�PDB�����)�
mc:cpmi�dbg��:�/  +����p�U   U��m�n3� X��d�~��~�a�{C�e����{g�+/�		^|f/s/i�u/~�
DEF �(�K�)�b buf.txt�/�/��W_MC�����Qd,53����ʇ>�Cz  B�p��B�Z�B�X��B��~B����B�<�C3���
q�Dv��D:��"Df��DR�t�DStD��a��=F�pgF�=C�Fi�WF��EF�2?F'jI�	ބ	6�����4���R(D~�2�/��ʄr3@à1/  TB��D�V@a  E�I�5� F*�� F�G$ˀF�[� GR�kNG�l��G��G���&H��G?֓�H��߃]���  >�33 G�ށ�x��@߂5Y�Ed��A���=L��<#�
 ��_�*~2RSMOFS���.^�9T1��D�E ��l 
� Q�;�P  x0_*_>TEST�")__��R���#o�^6C@A�KY���Qo2I��B�0��� �C�qeT�pFPROG %�(S�o�gI�qRu�����dKEY_TBL�  6��y� �	�
�� !�"#$%&'()�*+,-./01���:;<=>?@�ABC� GHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~�����������������������������������������������������������������������������q��͓���������������������������������耇���������������������9�Eъ`LCK�l��<�`�`STAT�c�_AUTO_DO���O�INDTO_ENB;���R�Q�Y�K�T2����STqO�~��TRL�`�LETE�ފ_�SCREEN �jkcsc� 	�UπMME�NU 1i  <�l�ol� K�u���FS����柽� ϟ���R�)�;�a� ��q���Я�����ݯ ��N�%�7���[�m� ������ɿ�ٿ�8� �!�n�E�W�}϶ύ� ��������"����1� j�A�Sߠ�w߉��߭� ��������T�+�=� ��a�s������� ����>��'�M���]� o��������������:#p)+�_M�ANUALӏ��DwBCOu�RIG��$�DBNUMLI�M�,1e
�P�XWORK 1k�_-<_N`�r�TB_� � m��Y0�_AWWAY��1G�@rb=�P�_AL� =���YҀ��`��_�  1!�[ 	,Q :&d2/o/��&�Mt�IZP�@|P�#ONTIM��d��&�
��e#MOTNEN�D�o$RECOR/D 1'kU2)?�!�O�?1-?&k� k?}?�?�?88�?�??? �?c?O*O<O�?�?rO �?�OO�O�O�O�O�O _�O8_�O\_n_�_�_ _�_%_�_I_�_o"o 4o�_Xo�_|o�_�o�o �o�oEo�oio�oB Tfx�o��/ �����>�)�7� t�� pu�����-�� ͏ۏ�����N�`�Ϗ ��o����)�;��� ���8���\�˟ݟ�� ��;�Q�گI���m���4�F�X��TOL�ERENC�B��	"�L�Ͱ CS_CFG ( +�x'dMC:\���L%04d.C�SVY� cֿx#A� ��CH�z �_/x.�G��},��R�C_OUT )�- z/��SGN� *��"��#��08-JU�N-25 13:�52��27�-MAY��4:3�8�]� Z��t�����x.����p�a�m��PJ�P��k�VERS�ION ���V2.0.11�~+EFLOGIC� 1+� 	�d��ٓ��p�PROG_ENB�\2��ULS�' ��p�_WRSTJ�N� ��"�EMO�_OPT_SL �?	�]�
 	�R575x#?�7�4D�6E�7E�50i�d�o�2E�d��j�>"�TO  .��l��k�V_� EX��d�% �PATHw A��A\��M�_�~+ICT�F��, '�`��eg��}�ST?BF_TTS�(�	���Eм`���� M�AU��ߧ"MSW��- )��},t���.�!��]l�R��v�����4SBL_FAULy��/��#GPMSyK�ߧ"TDIA���0����`���!�1234567G890xS�l�P�� ����//%/7/ I/[/m//�/�/�/�/h�/L0PV ���/�2?X? j?|?�?�?�?�?�?�? �?OO0OBOTOfO8<�x�UMP$�I� �ATR>�O�@�PME���OY_T�EMP��È�3p��4��DUNI	��w�YN_BRK �1��x�EMGDI_STA	��_��LPNC2_SCR 27[��_�_ �_�_�&�_�_o o2or�nSUQ13y_+?|o@�o�o�olRTd47[�Q��o�o���_ >Pbt���� �����(�:�L� ^�p������� ?Ǐُ �0�,p��+�=�O� a�s���������͟ߟ ���'�9�K�]�o� ��������ɯ���� �#�5�G�Y�k�}��� ����ſ׿����� 1�C�U�g�yϋϝ�ׯ ��������	��-�?� Q�c�u߇ߙ߽߫��� ������)�;�M�_� q��ϧ�������� ��%�7�I�[�m�� �������������� !3EW��{�� �����/ ASew���� ���//+/=/w a/s/�/�/�/�/�/�/ �/??'?9?K?]?o? �?�?�?�?�?�?�?�? OK/5OGOYOkO}O�O �O�O�O�O�O�O__ 1_C_U_g_y_�_�_�_��gETMODE �15'Efa �t|�_GgRR�OR_PROG %�Z%���Hog�TABLE  ��[1O�o�o�o�ZR�RSEV_NUM� �R  ���Q�`a_AUT�O_ENB  �u�SZd_NO�a �6�[�Q�b W *�6p�6p�6p	�6p�`+5pOastHIS�cXa�P{_ALM 17�[� ���6|6`+t���&�8�J�rx_�bp  �[�4q�R���PTCP_VER !�Z�!6oZ�$EXTL�OG_REQ�v9�y�SIZ�܄�TOL  XaD�z�r�A ܄_BWDo�%��fQ���w_DI?� 8'E�t�TXa b[�S�TEPg�y��P��O/P_DO�v$v`�FEATURE �9'EQ��Q�Handlin�gTool � �DER En�glish Di�ctionary��7 (RA�A Vis"� M�aster����
TE0�nalo�g I/O��p�1
0�uto �Software Updateb�� "/�k�mati�c Backup~
�d
!���ground E�ditB�  25�LCame�raT�FX� "L�o��ellT��Lw, P��omm9��shۡ�h600���cou���uct���p�pane� �DIF���tyl�e selectvѡ- /�Con��~9�onitor���Hd�tr�Re�liabT�ϣ(R�-Diagn�os��Q�	�H�Du�al Check� Safety �UIFc�Enha�nced Rob� Serv��q ��v	ԸUse�r Fr���T_�i�xt. DI[O f�fi�� )��\�endܰEr�ru�L��  pr$נ*�rO�� @����ENFCTN_ Menuİv��.fd`�TP �In?�faco� � 
E�G��p;�k/ Excذg�C���High-Sp�eܰSki��  �Par+�H���m�munic��on�s��\ap��ur�f�?�X�t\h8yU���connZ��2Т !�Incr��str)�8���M-6�KARE�L Cmd. L���ua��}��B�R�un-Ti�En�v�(<�@�I�<�+���s��S/W�"�H�Licen3se���� ad����ogBook(S�y>�m)	���"�MACROs,~��/Offse\��f����H�!�Y�M�1�MechStop ProtZ��3� 5
�Mi�4�Shif\��B;6S�MixܰQ�����H�Mode �SwitchY�M�ok���.�� ��MTt�Q�g�� �5��?ulti-T����ܖ�)�Posj�Re�gi>���  ! ��PA�t Fun<1��6iB/��R��Num�Y�3�G�P�/��� Adju<��	�/2HS�)�� o(�8�tatu����AD ��RD�Mޱot�scove&� #e�v������uest 867.��o�\���?SNPX b��Y�<��)�Libr%�
�Ort I���� "����.S�o� ��s� in VCCM,����� j������㣀/I�� 7�10�TMILI�BX����g�Ac�c����C/2�T�PTX�� �Tel�n��Y@����K�P�CUnexc�eptܰmotn¾� ������\m725����w�|5���  h640SP CSXC��i � j*�� RI�N��We���50�,��vrl�زmcen" ��fiP-��a���P��Gri�d{�play F� O/��? ��EL�R;�|�20��O{RDK�sciiw�oload�41d�;st�Patd���CycT�h���or�iɰ:�7c DatMa� qu6�2�0��*�������FRL�amc�K�HMI De��(����k��PC�φ�Pass�word�644���Sp�����D#Y�ELLOW BO��	?1�Arc%�v�isu����#ti�O�p�^�! 2��a6O�po�� t��ֶcT1o�����HT���xy�	�  5 $�t۠ig��1�0Ơ 41\+�J�PN ARCPSOU PR+�8b!�OL0Sup�2fil� �!��E@-�;�7croc�82��v����$ 12jSS�0e4�tex-� �I�7�So��tf�ssag�� e��У�qP��,��� "Tc �Virt��v�!�����dpn�
�J�3�SHADf0M�OVE T�MO�S O TԠ�get_var ?fails l�>P�U~1E���� Hold Bus %��h��VIS UP�DATE IRTORCHMA A�|{�vYWELDTV �S ]�DtS: R�741��ouiPb�}�y��BACKG�ROUND ED�IT "RC$REP�TCD CAN �CRASH FR�VR 62z1�SC�ra��s 2-D���r ) "��$�FNO NOT {RE��RED �`� m ��JO� �QUICKaPOP� FLEN m4�1S�Loc��gRT�IMQ%�#�FPL�N: FG��pl �m�r`�MD DE�VICE ASS�ERT WIT gPCV;PB�AN#a�ACCESS Mo .pc��Jo���Qui±�Kbld�mgUSB$ ��t� & remov� Pg�SMB �NUL� ;a|�FI�X��C��ACHI�N,QOL�`MO �OPT ՠa��P�POST0�WDUs C�wQAdd�`�ad���0io�2֫�$P�`W\0.$�0`O�IN&�P:�fix CPMO�-046 isskueC�J/aO-�0n�r130Т- ���vRSET VAR?IABLES-P{�ޯR3D m��vi/ew d��M��&��ea���b��of� FD�5P:N@x� OS-1y0`�h� sc���t��s ft�lo��7 WA�P�Z�3 CNT0 1T�/"�ImR�)��ca �Pu��PO�T:Whenape=wB�STY E�{1�t��ptKQdo /GET_�p �p��VMGR LOl�REAd0C~QW�~1��(�l�s�gD�EC�TpLpING /IMPR�DR(p+P�B�PROGRAM��ERIPE:ST�ARTU� AIN�-;�ӠM/ASC�IIzPÂOF L�q�DPTTB: �N�pML$me hP���`:x�mo&��allW`!�ӤTo�rc�A�U�HC�i�LpԸth�`n�@ �ch��/GEA�!�t�ou͐�RCal���k�Sign`� �ND�ԗThresh123��`��09p� : MSG_P�+0er  �Q�=Aܠzeron���0 H85��RI�mA�n�2D��rc:�0I��OMEa`�p�ONaP5�  נS�REG:FF-Д� �]�'���KANJI*��n��J��c�0as�n d�!OA im�mc �INISI�TALIZATI����~1wem�����dr+� LB A|�UWqminim�rec[�c!�R���}m$�ro -1>��S�ܰir��@ұJ�*1pdETw�� 5`?��I�ow u��< s_e 1lc��YbPM���p�Q���R`vR�&�lu\�3�Re �0�4q�q1#���m9 <a�arn���~��Box fo���*PRWRI�PW�S���v�09 F�pu�p�de-rel2 d�p� j��`━�betwe��IN�D Q���igE osnap|�us��spo TME��7TPD#�DO�p#a�HANDL 1\�k�`vR��ȀD�n�y�S�v�Yoper�abil� �T*�:� H � l\p��V�q�b�R�< p�a*�c&2O�`FA,�.�-QV7. f.v��[GT�pi�s���� ɠtmLin�e-Remark� �� RM-�` �W�#SPATH S�A+PLOOS U�IFc�+5f fig��pGLA����Vrp�������U�0the�r�V� TracD���tW�\b�s7���d�t�� n�@ I ���3:���dK�=y��it k8�d�wPayR![2]��^�1: g��s���dow�XQ��0I�S�q�qEMCHK EXCE C����MF +�Xah>�� 35\k��)���QBt���'b�d��[�c���e �`xk�S�� BUGrt��cD$`PETpȵ��f�c4��0XP�ANSI��DIG���@OoPmetTC�CRG EN��C�EMENT�A M�̀K {�`H G?UNCHG �`� �EXT�P�2�bQS��93 wP8�x�O�RYLEAKq � H5gyq�PLC WRDN R �sO /u�QSPE=p��G*�V ��$��tn720\3pGR�I��A�rT�PM�C ETH��pSyU7p�`  j5/^n�PENS�PN,���*P ont�`B�ROW�`!sRMVo ADDz CN �qDC���PT3 �ALA2@ ���pS�VGN EARLqY�R��ŰH57�GaJLAYҀEk (@M�PPD�p:*@H�S I`P��OUCH8���V�F�q�comH�x ���ERROR� DE� nJ��RO�C�URS8pI��Nx4q�-158n7��RSR xP#aU�p���Rqy�T�F�z�;�pk��t�� �gՂ�B�SY �RUNN�  a|�`�BRKCT�!�RO�p3@ \ap�SТ�AXxP���h�8+ q��ISSU�r} sPX�PTSI��K1M10_�I�PSAFETY Ck�ECK[��Á ������<#X�� ��TWD2�@�@�I{NV��D ZOp�5X��t�DUA=Ly� "M6�0�J"rF#�E��dPd?NDEX F�,t*UF�"Pʀ��0sFRVO117� A�PT6�KtqF�ALPTP247�7D6_�P�!;HI�G� CC�t;SNPX� MM��tq�d~�Vq�q#�
"��>DETEC�Tq*@RRU�qA�P�5p�9 y�)<9���7T��Pds� k�	���!Q���� t\4A�;A0�o2 "Ke@" 8@�HI�qXF8@4@H�PRDC"�
�aMB8@�IXF�b���zOX@8@����a�G}E�B�Ccs�cr�J8@�Ndctrld.�A�NZE�A�5��Q��!�`�Df�8@�`m�878�Q-z;� ��� rm`�i
��PR̠78�@�RI8@0q�Q ( ~\Mp��0t��!{B8@�\tQ<OX�St0�32hB3nO�Vtp�A�@gLCF�L��� �Rplcf���J8@�WTamai�E8@mubov2_miTA�O�S8@�U`T[tT�AqPr67�4xSShape GGen��8@j�I�[R�`�@8@T����%qc (u8@��II�^��Q~C�a�[8@;Ynrsug0�4� � 4�C�tMr68@�r5hB5��zVnretsp e"r�Po�wng0bGCRE�Ka�ޠ��DAT�E�k�creat.�q�M��a�oksqgtpa�d1P��(�tput�Zj�{�������܆2�8@����Q����sl�o��� �hex�H�TB�8�ď�ke1yH�8@�pmZb�NbR�u7A+�nrgc8@ UQ�pp�bUZ�dp0a�j921xSpl.Collأcq�\A�b�RNq�UA� (J�8@ip�_�WA��_�Y���a7hB7�ͦt�p[� "TCLSx9oKb��clskyht[��s�pkckZd ���$�TQ���dA�r�x�710a- KA�REL Use {Sp�FCTN9��a�7l�0s0a�� ( ���a��~C8@��MI���c8hB8"   ��8@ v	��v	   �lmatea99�qM����E�mcc;lm5�CLM;�� ��j��E�et���aL1M	�h�yasp,���?mc_mot�B�N���8@H����Q��su�'��Q�ȕ�䅮���j�oi#�ߕ��A_l�og�Z���trc�B����ve�ϓ�v���QWX��6�find�erxSCente�r F1�lSw52a0��ha6rX� (<�cr,�Q�Ձfi�Q  �NH0�I�ۡ���A8@�uL��tq�a "F�NDRVϳ���et�guid�UID �C8@���������TA@�nuf;��P�����C�B��_z�Ӡo��qG������l���f�ndrTY��2䁴t�cp"�,qCP MtF�}38@517��6s38�E��gf6 ��(��K��Q��-�X�L�A�tm6�P�� ���Q���	�����tm�Ĵ�b8@aej��TAiex���aP�Aa�ذ�cpr�m�A��l�_vars��
��dwc7 `TS��/�6��ma7A�F�Group| s�k Exchan�gJ 8@�VMASK� H5�0H593� H0aH5@� 6V� 58�!9�!8\J�!4�!2���"(�/���;OMI� `@a0�hB0�ՁU4U1#SAK(x2�Q�0I�h�ӂ)�mq�bWzR�D�isplayIm�Q@vJ40�Q8aJ�!(P��;� 0a���0��� 40;�q�vl "DQVL�D쌞�qvBXa`�uG�Hq�OsC��avrdqq�O�xEsim�K�40sJst]��uDd X@TRgOyB�Bv40)��wA~���E�Easy� Normal Util(in��K�11 J553m�0b2v�Q(lV40xU�)��������k986#8Uϕ�|�rP "NOR��dw d.a}oKksu�O�W����OY�W`�j0�6�H� �menuuyP6�Mx�`wRX�R577V��90 �RJ989F}�49b\�`(�fity�����e��<?��Vsmh`��8@��C0�Sv�q�8����w�pn "MHMN<��ޣx�Ay`�o��3�u�`f�І�x�t ��tRzQ��LV��vP�#tm���|I�1{oPx" �2|���I�3I/B��odstǏًmnx����}ensu_�	L<���h!!��Rt~��huserp��0Ҹ�ʐcM�_l�xP�oe��рpoper�����xdetbo /�l>�x���Ps$p��`���OPydspw�eb͓��z'R��u�Rr101&S՟{tb�`2�Z4�30������`4�
�4�5���KQ�m[T��dUCalG40`�Q)p40}������9;��DA��? v	LATA�umpd�\bbk7968��68c�f�bl�41969y�9и|�D���bd� "�BBOXêM��s�ched����m�s�etuM:�����ff���40��n�41��8��40q�col��|��1�xc�ؘ���li ��X�0���j��&�8��4 <�ro5�TP �E�#��ryK412r��;�(T+Q �Rec'�ʈ1Iw��84�����Ak97�1��71�;���p?arecjo��Q�NS�[T���dXra{il| nagek��M ,QT2 *� !(�ĜR%<x�80P!bh��p��4���4�yDgl�paxrmr "XRM�g�l�brf{���n���kl��9turb�sp��㧑- �l0s15	�g�625C� Mh�+���)89��	+��B6��o�ҹ��x�7�q40�����pd "TSPDx�=��tsgl��l�:dQ���8Bc1t���K�vrE�a�ܮ�����  ��!���21��`( AAVM� �2�0 �@fd� TUP him� (J545� l)�`8 616� %�VCAM� ��CLIO] (�0:�5& � (F\ MSC ��Rt"PBsSTsYL�D!28 :2�\ NRE F2h S�CH6pDC�SU tpsh ORSR �r�D!04�SEI�OC& \fxh 542 LEX"� ESETn�8!H ���sh8 7H �OMASK�Ø"7>�.�OCO*`x�!0�3"6�!/400:66�$ G639.6[8LC�H!6OPLGR70=3
5MHCR��0�C� (! �06�A.�f8!54
��00D;SWb 588�180� �h!37 88 K(D�"02C24��N�27 q9�25���2-6�05��9�PRST bB/FRDMES�!zB��930 _ N�BA  6� HL�B 3 (~!SMވ@ Con� SPgVC �8!20z���TCP ara�m\TMIL� A��@PACET�PTX �@p T?ELN 96��2�9�%UECK��r� UFRM et��P!OR ORP I{PL%CSXC�0�j�1CVVF l� FQHTTP �stA")�I#� CG�HP8ZIGU�I�0�hPPGS oTool� H8�@�djZ��!@�h!6�3�%�@32Q\�31� B�h!96�%R6�51�Rs�!53 oTFAD�R41��8"1 ��oo�"9:��41775�"/@�P�VCTO�@�U�!�sh!80�%PRXyY�R�!770 �b~8 885 ol3P2� L� аdi� �`�ڳh LCP{Q� T'SS �b�26:���^�@CPE �HT@�VRC~�tQNLy ��@002 %�b	0dis� �`7� <��a\0�T�`1 ��`en�b4 6582�`)FU02Q0Π�o`p�Ptu�r4 d$r5N��RU0p@�nse�QJp1 A�PFI[ Jp3�g3}4�g40 al�xrE1t44w466� ts U0  7v��0O��r5�e�p7 �p "sw�a61d:��r4��r5 Qp!wGr`�$�p8R�"s�P`tQ�b�36w717�w8`�v83���r�8�&:��pOq8�8 _"rkey8�9F�v�a90�91 p�p#@��� �D095�g[97*pur�A1@ d���P|P�q1�0QplSq1p#4��]a!sM1@sl༂8��H��\1�d1�`��v��@{�14p�ae��5# h2��`�6ޣ��7�f1p@��d�YpCq(d�ـd�1�`uq���� Cu1< Oq� ��7&ReU1$ �u1�Pϱ�� ��@- WQ1�58 ase C渒9 B��60 �82ń�p���4 (Wai��`吢!���7E��8�EU1&P`ro9�<�1��<�2��<�	0��T��"l�5J�l��cC���9%�MCR��P��2�`�Q2@96I7�Q��8��9Z�A2TPB���P�2P7�U5@�o���
�58�`U���3 w����?A�E�1��c�qAw�l��A�1��512# f��1�u5Р��"�a5p$��56�+aĈ�Q5h��Ұ�1 �@��pp�b[�538 xaB��|p�4Ⱅ2�11/q5�p�4U=5�P16 (߲�P z��0��8�P��H���p�e5`�e5(�/�P`bbf>�X��$�Z�U�5d�\�� X�7 	  ~��8 k_kv���79 s�82 &�H5��E6���p�����h���ñ���3�J"�`��4 3Ȥ5�9ѧ6�0t���8Ⲗ6D0$�$�4 7���!���<�j67?0\tchk<�P`s��<�B<�90���7�<���<�\K�<�q �Ӻ�A�C<���q�<д��<�t��sg<�lIc���FA<�H���<���<Я���<�hk ��<Щ�B<е�o�<����<��K�<�dflar��<Ш��� ��@o�`���D�;�<�gEvam����B<гoќ���<а�KЀ�creexl����P�`��<���|���j6<�=s��prs.`��� \���<�7������fsgn��P�b�t�at��<�L��1|B !�svsch/ � �Servo S΋�ule>�SVS��44�1u�_<���� (����ched��,��~��A\�� �� B���B�qA�h���cj�� � 5�1<���Ә�p��css "ACS <�&(��6� ������c el���Q�����torchm�s�<�- T�Ma�`Ѵ���09 J5�;598 J681s�7� 8��b���<Чa����te,s�����/�E��� m��ARC..�� 1q�4�!=�,�C�tc�pA�@t����f� F����7#�2x�SE�r����UtmS�09610'���RC�������� p��96`G= '��"H5W�@���L���\f� � �PATb���`!a4U�#!Stmt��E ��� �pM�A�!p��z�2?�i�n_<�X��r�X e/cW����V����etdl�vߏ\oveto���܏���mmonitr`�\��|#�0st��?.6a��PP�����! Q�!y`�`asme �Arol�6c�43�0 �pl���01� 25��  �<� v	�v	�A>@�818\n; <�s�I�B�2�pMPT�P"��C�1mocol��,��CT�v�'!`� �A���8P53��y`Touchs�s0�`��<��J5��@�Ѩ`mP����n[P Q�a,�E�a��IPL&
�Pth�A<�KF#xR�m;�Qetth�THSR'�q-�Rt���o "PGIO��#!$s�ISwka�"cWK��!�MHqWH54��5w5n/"�Sm/��@ 7�*�da��8`!w/Ac��tsnf Tk�/�#@gb�a��u`��^m�`Au��Zӭ�ܱQp��@��#���Ka<��M��t5QtZ�a<��d�FS5GK����G�1o1r��dW��64��tP@x���P ����x,� �?$���P<�Z4e�7�g "SVGN�.ox�copy "CO;�Wj$�O�A�9� "FSG�ѧ�%�7��_��f� wQS�WF*!"(�sgat�uɀ���_
��tpN_TPDo��9�79�#dߎ?���h��GAT���!#��  �Гf�` �@�"/� �w�Z� �b?6 ?� ����� ���E �8��M� �chrT� �K6K� �sms� �o6��ѐ�gtdmen�?3 �?��� ���mkpdtd2 ���, ���pdQ�X� ������ ���mvbkup�. �[�C�С��mk3uno��prp���Gmkl �4��s ��niU��� �ldv9rw���glg�4��� ��棑��aut7�.pб�旐 �ַ������su3� ��@�� �Ƿ� ���\ �6�b2X� ��&�� �x����A4�  ���B   946�" ��fB� �t\p�aic\p4k947 ���F#���� ��ictas���pa`���cc:�<��8o�����gen�� �I ��F�lnp � �Ď��stf@��1��wbO�c��Ջ�`��߄�vri�ߢ�а�-T� ���p�flo�w� OPAc��ow���R50qtS �#T� (A��4�#�0��pѣV�cu3�Q0F� ��SI�ac�����46����s&��p�a��!!���� ���55�b �o)�p���0�|��
�afcal3�P� ��f��}���`�f��m	߳�p�d�m�/���a/��$C`ѷ��� �! trac�k\P� 0�ine/Rail Tr��]TJ�69W�T  (L��8(`љT.�`� %��D��P0� (��8�48��_ɛ�₇�4����� �3b�b3���alV@ �NTf���%��I�in]0m���aen������&?5�8c@Itst3@�� $����`�,R9�%����0氱%��po�peners-OW dDev��F�M�6W���|A�Pc"�l!esv� �,��R�V$�Q���U<�V$ �k)9j �6��# ��ȼ��%paop/!O�PNU�V ��2c#elL��8g_��8/�6��tscG��$Ѐ�V!�3� 5vrCop�ߡ�7`�n( `�V"2D�a V'O$�:S9��� Pump E��jQ�@�" ��!
��@бMSC#�@��)P���AC�`��� � �v���� \mh/plug�@g�"�7P��uK")㠱io�7�CJ0��E�LI�O q1g 7A93շ�5 q9 t����]4rb ST��R�ÞCPJ989�P�L�SE�' �e C3Q(P �/Ov���o�P� ? I1�R����55��f�I1`�tcwmio��MIO������Utco1"CL�01V �cBK`iEo��uM?���Sl� I0�ߢ�Eg �o���fb �tI4\onfdtI����e%�p27�Inste�TB CoMIoo1E�R�(do554 (;r>Ex�,��nR##ipc��/>��qp5���
@oQé�1�p����7/o����ra�pd�CD V_��rP�֮��qp2Gcnd��s �p��a�o�r`҄�S��"�bc�a�c���2kI�<�?A�pcrt���or0�qd#��"���3p�+���D��Џ��vr2k�0���AG�.�+��cho�;�u�C��(� �uV630 �fwe P�mී�@�X��`��TX�� ��>d�chp "_��(	�3�����8����\p3�v�������9�3�1 ������low�[ͧ���c!hk���㳦s��s?Ө0�i�1h���2�� i�w����s?1*�`-	�:�O��vr�������0�'���PFR�APWat?1rn�eE�P�sp�& ac5�� _A�rbo#�, �a��g�������z�Qs<�ICSP+� 9_����� ��F�A9PH51�IQ93 7��HX6�hQ]PVR`S5��fPR�6 iQWPR� (�P!am S�u�"�A�I0�tppr�g�0���`h�@2atk932�!��E��^��asc "8�C8��S>i�atp�"��d�@1I�
g�ds�blfltJA�Qs�able Fau�P{C!��EV0ex~/!DSB (DC��t�$�p��X 7�@� �� 5��Q�t3*��~���td9� "`!%�(5��sb9������\	�6#���@�5�p$D@550-A�djust Po'intO"tVJ�Rs�z�䐄��!�X_�Yj���0\sg��4x��}7y�\ada�O"ADJ���j�Q�etsha<�SH�AP�sŭ'jpo �r4�t�!��$ �(�C|�	Tk!bRP�KAR/Qiagn/ostì!O!vV66 J`ew0��(�L���/�&krlde� ��PP�� �hU b���r3�Pyp?q��DBG2C��� �X�o�1U��� ��WT`�@i�pJCM�aipper Opv`1Se}�78 (MH G F� ;":�&##�� a��x�֕$��388�C�����#��9.�9�C��g##PPk�Q��8 �!�_"$�"��=0%�P� �A $��_�#%0AQ�C�~2 Mat.HandlE��!= &�pq MPLGET�0�1(�3�Tt&P�Sٰ' �B�1��B0����&p� �H��PP �'p��@�C 7PP	�TG�tD5�}�m�q�Afhnd �"F_R  ������PP	   pxT?Q���P(Pa���To�����?�p�mpaO��JP ak925��2`@O�JR	psQ`B2�unLHP�T7gse�GSo1�O�W�QT��v !�R��Ptp~���JRdm�on.�@��V�!ns�hYvr�QJ�g�Q`�o�jY�HS~7sl�f] ��pen�PDnRp(R&���ɐ823'� �ٔq���g� ����� 1�� S�� ? �c\sltQ�!|QE�P��a �rtPg��P�� �v��"SEDG8�s0.�qtdgY T�� ��vP`ho�s`<` ����qc�`g
�e`� o�w�a@o"�ile6�H�e�ȅnR��� �e! j517�>Ճ��J%��e�`��Q4��Q&�!L�!F�J�=�o�5�z/l17���_�œ���`C0C�  ���LA/NG j��A��p������gad����#�jp�.`��4�Ē�ib�0��s�Ƒpa����&���j539.�f�,Ru� Env
�����2�3H�z�J9������h�Ф
Ҕ���2��2���� (K>L�n-TimФ������p�3�TS�����\kl�UTIL�"o���x�r "QMGl��!������1 "��S�T3�\kcmno��SФ�T2���ut�.�l�readc�}�exPY�ܤ�r��\��l�҄Фw�3��2C�*� -�C�D�E!Ĥ� .�4�C� R CV̴�҆��\p�Р���p�tbox��.�@��cycsL�:�RB�TE�veriOPTNE���;ӕӂk�e�ߦ�a�ߦ�h�g�ߥ�DPN��g�p.v��r�ptlit��0�4��te\cy���>�tmnu3`�r�����5UPDT�������駣���ite �� sw�to�,���oolB�F"�Y���Q��(q��gr3��䪒���"�䴁w������߳��s��������������lS���bx A"O�� ����l��`��P���A�l\t��� ��������	�Co�l�e!��R C ��r��&r �m;`��Chang�Lq�T1 �rcm3�"��
� 6���"����sPa7���"��22B2��2D4�57�� CC�FM�H��accda��Q�c' ��KÕ0���K!����m o!���,$Á��! "
����/�/����	�Y�,$��)�,$sk(����m rC%tS1,$�+��k1�%unc.�,$oñ�1��sub������1��cce �5/!&��-/?-W/i&vs�}/�%#�#�/��.C��/� C%
�@?  U �&+��F:qt�
pD�Ѓ D	 � U�:7�Dxmov.�P��DPvc\5Q�tfr@PeC_~UYgeobdtg_y[tu���P���PTUIt�P�Sx�_�^z�_��\var�_�\xy\�_�[pcl`c�P脆�P�Ue�Pgri�psuaoskuti����ovfinfpo}��o�j�b�P���Qud\�aX��Pc�\Rrp�Qnƅ�P�v�P)t�m#qƆ�P�v�a+ro�g�a��\Q�?a+rp#al?a{�{spa��@�P�u�Q�t�_TZp�0<�osipkag3r�o>vlclay(�:�t�pT�d�pu?a�c�A������KtKa�P䒏��qTf|rdm��{rin#r���As� �2���|s�PLd�v�tv��v�h�0��ystn* џ�y%t'�1�p��D�p�uϑ#�ul�@o�W6�92�siupdl�]�Fo�vr�on��`1L��z�`\�r���il3�$|l4��ǉ#q5 4FyB�Տg{�`���{�wcmס���wxf�er�UYtlk2�pp߿UYconv��sicnv�Qʯx�ag��H�Z�lct�`ao�=�p��׭nit0믁�3�������  �� ?v	�v	$��alϑpm�r&�B�eWa���f�%�� ����I��߬�u�ͬ�KamT�f���c��w��roǁ#�5�����?� sm��y�a��y� ��������`����͐ϑ��p��m�Wa� 1���A�6�S�e�X� �ψ�\Q}��������� ��ĥw߉�西߭�� �߮�#q0��rs�ew����1�a��z긱n�@�.�۲;�d�������  � �Ad	T$�1 �p! P��e �Ne 	lf@C��@�s/�  ?�����8�� �������r�eg.�C=��o�99 ~@�����$FEAT_�INDEX  �z ���e� ILECO�MP :��=�1!!z�$#SETUP2 �;1%;"��  N f!$#_A�P2BCK 1<~1)  �)��/�/  %�/�/e4 �/�/>%�/$?�/ H?�/U?~??�?1?�? �?g?�?�? O2O�?VO �?zO�OO�O?O�OcO �O
_�O._�OR_d_�O �__�_�_M_�_q_o o�_<o�_`o�_mo�o %o�oIo�o�oo�o 8J�on�o��3 �W�{�"��F� �j�|����/�ď֏ e������0���T�� x������=�ҟa��� ���,���P�b�񟆯 �����K��o���� �:�ɯ^�����#� ��G�ܿ�}�ϡ�6� H�׿l�����ϝ���t@)t Px/ 2� *.VR��߅�*�@߂�F�j�T���PCrߛ߅�F'R6:����V���z�T �!���K�� ��q�S�*.F�ߢ��	�Ӑ���x^����STM ��'���S����iPendant? PanelS���HI���9���U�������GIF0;�p�������JPG���;��]oR�
�ARGNAME.SDTy�>�\"����Rc	P�ANEL1Y�%�>��e�w��2 �A/�//���/�3_/�/��/p/�/?�4�/I?�7?�/?��?TPEINS�.XML�?>:\��?t?�1Custo�m Toolba�r�?Q�PASS�WORDg?w�F�RS:\:O�? %�Passwor�d Config {OR��OSO�O�O��_ �OB_T_�Ox__�_�_ =_�_a_�_�_�_,o�_ Po�_Io�oo�o9o�o �ooo�o(:�o^ �o�#�G�k ���6��Z�l�� �����ƏU��y�� ����D�ӏh���a��� -�Q��������� @�R��v����)�;� Я_������*���N� ݯr������7�̿޿ m�ϑ�&ϵ�ǿ\�� ���y϶�E���i��� ߟ�4���X�j��ώ� ߲�A�S���w��� �B���f��ߊ��+� ��O���������>� ����t����'����� ]�����(��L�� p��5�Yk  �$�Z�~ ��C�g�/ �2/�V/���// �/?/�/�/u/
?�/.? @?�/d?�/�?�?)?�? M?�?q?�?O�?<O�? 5OrOO�O%O�O�O[O �OO_&_�OJ_�On_ �O_�_3_�_W_�_�_ �_"o�_FoXo�_|oo��o�o�`�$FIL�E_DGBCK �1<���`��� ( ��)
SUMMA�RY.DG�obl�MD:�o*n`�Diag Sum�mary+8j
C?ONSLOG �qn�=qCon�sole log��7kpMEMCHECK��2���qMemory� Data3�;g�� {)�HAD�OW(�����C��Shadow C?hanges���c�-��)	FTAP�����=��q�mment TB�D;�;g0<�)�ETHERNET�0�`n�q~���=qE�thernet ��pfigurat�ion��B`%�DCSVRF/��'�@��C�%� ve�rify all�C��c1p� �DIFF8��0�ůD��%Z�diffǯ{��q�1�������J� X�q�|�=	�CHGD�&�8�ͿD�ܯ������2Ŀ����R� `�yτ�GD�.�@����D�����FY�3�ϳ���Z� hρߌ�GD$�6�H����D�����UPDATES.$��
�ckFRS:\�"�c�>qUpda�tes List�c�`{PSRBWLOD.CM��blN����e��pPS_ROBOWEL\�6o+� =�loa��o����&��� J���n�����9�� Jo���"��X �|#�G�k �d�0�T�� �/�C/U/�y// �/�/>/�/b/�/�/�/ -?�/Q?�/b?�??�? :?�?�?p?O�?)O;O �?_O�?�OO|O�OHO �OlO�O_�O7_�O[_ m_�O�_ _�_�_V_�_ z_o�_oEo�_io�_ zo�o.o�oRo�o�o�o �oAS�ow� *��`���+� �O��s������8� ͏ߏn����'��� � ]�쏁������F�۟ j������5�ğY�k� �������B����x������C�үg�v���$FILE_N�P�R]���Y�������M�DONLY 1<���U� 
 � �ۿ(���L��5��� Y��}Ϗ�ϳ�B��� ��x�ߜ�1�C���g� �ϋ�ߘ���P���t� 	���?���c�u�� ��(����^����� ��$�M���q� ����� 6���Z�����%�� I[���2�����VISBCK�����ų*.VD��*� FR:\�V� Vis�ion VD fileVd��� ����	/./�R/ �v/�//�/;/�/_/ q/?�/*?<?�/`?�/ �??�?�?I?�?m?O O�?8O�?\O�?�?�O !O�O�O�O�O{O_�O !_F_�Oj_�O�_�_/_��_S_�_w_�_o~�M�R_GRP 1=LeC4 w B�`	 ���lo~li`۬B���D��f�nӺMT� ��� ����e `i`a�o�khb�h�o�d�cic.N����L#�L
��+N���H�M�E��|��i`?{��Aǿ�@i=F
��A S�8�[�ol}A��A���A���s����p�l}F@ ��qhq�y�~g�fF�6�D�MqD��� BT��@���Ô~pD��6����l���5��5��|���~�� B���B�%A���B�>zBZw��~A�B*~�B6��A��9�B O7B�B0l叐�A��� ��A�܏e�P���t����@�bo=���@�	Ƙ� ���Ο��+��O� :�_���p�����e;BH` �Ă<��a?T#=����'�d
��Z��WZ�qW/�FX
��A@���@�33;@����\��[���ѿ��@��񿋯 �*��N�9�r�]ϖ����<�G�=��<�m]<��+=~�m<c�^��8eN7���7ѷ7��x7;��51�@��	ߤ��?߾d2^`UYb`�b`������F�`Үb` b`:�0�����C�^o �߂o�o�߸o��o��  ]�(߁�l����� ��������#��G�2� k�V�{����������� ����1 �� -�)����� ��0T?xc �������/ ')�'/M/_/q/8��/ �//�/�/�/�/?#? 
?G?2?k?V?�?z?�? �?�?�?�?O�?1OO UO@ORO�OvO�O�O�O �O��_��J����`_ *�_N�_�O�_�_�_ �_oo'oMo8oqo\o �o�o�o�o�o�o�o �o7"[Fjh �x�t��!�� E�0�B�{�f�����Ï ���ҏ����A�,� e�,/���������/� J����=�$�a�H� Z���������߯ʯ� ��9�$�]�H���l� ����ɿ��ƿ���#� �O�OV� _z�D_V_�� z_�Ϟ_���
�C� .�g�Rߋ�vߛ��߬� ����	���-��Q�<� N��r������� ���)��M�8�q�\� �������������� ��7"[Fk�| �|����֟3 �WBg�t�� ���/�///S/ >/w/b/�/�/�/�/�/ �/�/??=?(?:?s? :�LϦ?p��?�Ϧ� O ��$O��T?]OHOZO�O ~O�O�O�O�O�O�O_ 5_ _Y_D_}_h_�_�_ �_�_�_�_�_o��@o 
�go*owo�o�o�o�o �o�o	�o-*c N�r����� ��)�;�M���� �����ˏݏď�� %��I�4�F��j��� ��ǟ���֟��!�� E�0�i�T���x���ï �?�?��O��?OO �t�>O������ѿ�� ο��+��O�:�s� ^σϩϔ��ϸ����� � �9�$�6�o�6o�� Zo��R���������� 5� �Y�D�}�h��� �����������
�C� U��y�����d����� :�����+Q8 u`������ �;&_Jo ������// گ4/��x�j/4��/X� n/|��/��/�/!?? E?0?B?{?f?�?�?�? �?�?�?�?OOAO,O eOPO�OtO�O�O���O �O_�O+__O_:___ �_p_�_�_�_�_�_�_ o ooKo6oooZo�o Z��o�o�o�o��xo 
G2kR��� ������1�� .�g�R���v�����ӏ ���	��-��Q�/ */��N/��r/�/ޟ�/ ��/)�D�M�8�q�\� �����������گ� ��7�"�[�F�k���|� ����ٿĿ���O�O�O ��W�B�{�fϟϊ��� ����������A�,� e�P߉�t߆߿ߪ��� �o��+�=�a��� ��p���������� � �9�$�]�H���l� ��������������# G2W}h�p���$FNO �������
F0� ��  #�1 D|��� RM_CHK�TYP  � �\q�� �� ��{OM� _MIN� �m����  �X� SSB_C�FG >� ~�Jl��Aj|�TP_D�EF_OW  �m���IRCO�M� ��$GENOVRD_DOs����THR� d�d�_EN�B� �RAV�C_GRP 1?3� X�e/� �/�/�/�/�/�/�/�/ ? ?=?$?6?s?Z?�? ~?�?�?�?�?�?O'O OKO2OoO�OhO�O�O��O�O�O�O�ROUr? E� q�������8�?#�O__K_m_o_�?�  D3���_�E�_q�@A��\B�����R��>Y_6 SMT<#FC-�Ufoxo|�o�HOSTC,s1GY?��_k 	�h�k�o2�f�oyeC Ugy�z1�������p	ano?nymous�5� G�Y�k�w��o�o�o�� ����*�<�� `�r�������ˏ	�� ���&�8������� �������ȯگ��� M��4�F�X�j����� ݟ��Ŀֿ���I�[� m�ρ�fϵ��ϜϮ� ����}�����,�O� Pߟ�t߆ߘߪ߼�� �/�A�C�(�w�L�^� p����ϸ������� ���a�6�H�Z�l�~� ����������9�  2DV��z�� ����#��
. @������������ ���//g</N/ `/r/�/����/�/ �/?Qcu��/[? ��?�?�?�?�?)/�? O"O4OFOi?�/�/�O�O�O�O9m�aENT� 1H[ P!\^O_  `_ ?_._c_&_�_J_�_n_ �_�_�_o�_)o�_Mo oqo4o�oXojo�o�o �o�o�o7�om 0�T�x��� ��3��W��{�>� ��b���Տ������� ��A��e�(�:���^�𿟂�㟦�QUICC0�̟ޟ?��A1@��.����2���l�~�߯!ROU�TER௼�ί/�!?PCJOG0���!192.168.0.10	���GNAME !��J!ROBOT����NS_CFG �1G�I ��Auto-s�tarted/4FTP:?�Q?SO Bχ?f�xϊϜϮ��? �������+�߿�P� b�t߆ߘ�6��� ��(�J� �1�C�U�g� 6ߋ���������x� 	��-�?�Q�c� ?2? D?��������� )��M_q���� :���%t� ����m������ ����!/3/E/W/ z{//�/�/�/�/�/ 6HZ ?n/S?�w? �?�?�?�?�/�?�?O O<?=O�?aOsO�O�O �O�/
??.?0O_d? 9_K_]_o_�_PO�_�_ �_�_�O�_�_#o5oGo Yoko�O�O�O�O�_�o &_�o1Cog y����oT�� 	��-�|o�o�o�o� ���o��Ϗ���� )�;�M�_�q������๟˟ݟ�ÿT_ERR I������PDUSIZ  ��^���$�>~=�WRD ?޵�w��  guest+�}���࡯��ůׯ��SCD�_GROUP 2]J� �`�51��!��L_����  ��!�	 �i-	�E����Q�E EATSWILIBk�+���ST 4��@��1��L�F�RS:аTTP_AUTH 1K��<!iPendCan�������!KAREL:q*���	�KC��.�@��VISI?ON SET���u���!�ϣ������ ��	��P�'�9߆�]��o޽�CTRL �L��؃�
���FFF9E3���u���DEFA�ULT��FA�NUC Web �Server��
 ��e�w���j�|���������WR_CONFIG MY�X����I�DL_CPU_P5C���B�x�6�w�BH�MIN'���;�GNR_IO��K���"��NPT_SIM_DOl��v�TPMODN�TOLl� ��_P�RTY��6��OL_NK 1N�ذ �� 2DVh��_MASTEk�s��w�OñO_CFG���	UO����C�YCLE���_?ASG 1O��ձ
 j+=Oa s�������p//r�NUMJ�� �J�� IPCH��x��RTRY_�CN�n� ��SC?RN_UPDJ�����$� �� �P��A��/���$J�23_DSP_E�N~��p�� OB�PROC�#���	J�OG�1Q� �@��d8�?р +S? /?)3PO�SRE?y�KANJI_� Kl��3��#R�����5�?�5CL_LF�;"^/�0�EYLOGGINʦ q��K1$���$LANGUAGgE X�6��Y vA�LG�"S��V������x��i�j�@<𬄐'0u8������MC:�\RSCH\00�\��S@N_DISP T�t�w�K��I��LOC��-�D�zU�AzCOGBOOK U	L0��`d���d�d��PXY��_�_�_�_�_ nmh%i��	kU�Yr��UhozohS_BUFoF 1V��|o2s��o�R���oq��o �o#,YPb� ����������(�U��D/0DCS� Xu] =���"lao����ˏݏ�|3n�IO 1Y	G �/,����,� <�N�`�t��������� ̟ޟ���&�8�L� \�n���������ȯܯ��Ee�TM  [d�(�:�L�^�p� ��������ʿܿ� � �$�6�H�Z�l�~ϐ�8�ύd�SEV� ]]�TYP�$�`��)߄m�1RSK��!O�c�"FL 1Z�� ����߯���`������	�:�TP5@����A]NGN�AM�$�E��k�UP�S PGI|%�1�%�x�_LOAD0G� %Z%TE�QѼ��MAXUALRM;'�I(��~���#� V�#a��CQ[x�8��n��"�10�60\	 �F�	 �Ϣ�������������  D'9ze� ������� R=va��� �����*//N/ 9/r/�/g/�/�/�/�/ �/?�/&??J?\??? �?k?�?�?�?�?�?�? �?"O4OOXOCO|O_O qO�O�O�O�O�O_�O 0__T_7_I_�_u_�_ �_�_�_�_o�_,o���D_LDXDIS�Ac���MEMO�_AP]�E ?��
 �5i�o �o�o�o�o�o�o��ISC 1]�� �oTd��\n o������� ��I�4�m��f��� $���������!�� E�ƏT�f�:�����ß �����z��ܟA�,� e�w�^������~�� ���� �=���L�^� 2���������߿�r�� �Կ9�$�]�o�(t_MSTR ^��~��SCD 1_xm�W���S������� =�(�:�s�^ߗ߂߻� ��������� �9�$� ]�H��l������ ������#��G�2�W� }�h������������� ��
C.gR� v�����	� -Q<u`r� �����//'/ M/8/q/\/�/�/�/�/��/s�MKCFG �`���/��LT�ARM_2a��;2 �#\`|Y>G`METPUT`��"����NDS?P_CMNTs5086�5�� b���>��"1�?�4�5PO�SCF�7�>PR�PM�?�8PSTOoL 1c2}4@p<#�
aA�!aEqO G]OO�O�O�O�O�O _�O�OA_#_5_w_Y_�k_�_�_�_�_�Q�1S�ING_CHK � +O$MODA�Q73d
?�7:eD�EV 	��	�MC:MlHSIZ�Es0���eTAS�K %��%$1�23456789� �o�egTRIGw 1e�� l��3%��?   A$�ÜfYP�a,u���cEM_INF� 1f>7 �`)AT&�FV0E0N�})��qE0V1&A�3&B1&D2&�S0&C1S0=>�})ATZ�� �H�E��q9m��xAu���X�������� ������v� )���я��П������ �*��N�����7� I�[�̯ן���9�&� ��\����g����� i�ڿ������ï4�� XϏ�iώ�A���m��� ����߿�ѿB���� ϊߜ�O������ߟ� �����>�%�b�t�'� ��K�]�o߁����� (�_�L���p�+�����������.ONITO�R�0G ?ak  � 	EXEC�1�#234�5�`78
9�#��x xx*x6xB xNxZxfxr�x22�2�2��2�2�2�2��2�2�33�3aR_GRP_SV 1g�y��a(�Q>`�?��뿲���cj�?�ZF@gK�	Hm�a_Di���n�!PL_NAM�E !�5
 ��!Defaul�t Person�ality (f�rom FD) ��$RR2� 1h�)deX)dh�
!�1X d�/d/v/ �/�/�/�/�/�/�/? ?*?<?N?`?r?�?�?�?�?�?�82S/�?O  O2ODOVOhOzO�O�Ob<�?�O�O�O�O_ "_4_F_X_j_|_�_Lh�R� 1m)9`=\b0 �_pb��Q @D�  &�Q?��S�Q?`�Q�aAI�Ez � a@og;�	l~�R	 0`�4b@4c.a�P�Jd��Jd�Ki�K��J���J����J�4�J~���jEa�o-a�@�o�l[`@�z��b�f�@�S���a�Q�o�c�=�N���
������T;f��`���l[`�*  �p�  �$p> p��$p��o?p?�����	��o�Bntr�Q�s�kse�}�l�p��  �pu`j7  #p��vks��� 	'� �� �I� �  ���}�:�È6�È=����N��b@�^�d��n�Q���{�RȒx���nN. ��  �'���a�`@a��@�t�@p@�p@CpCR0�f0�+pB/pC3}=�P�@%�Ea�b�oo�$|m�����gA%���. ���z�`�P���QDe����˟��(��m��� �t O�� ru �4� �R�c��s�' :�u�a�P�`? �?�ffb�!������7� ���گ쬛af��>������iP�P;�e�S�xEa4f�u�>LX���s�b<	�I<�g�<#�
<2���<D��<���
vo��¯�S���S.���?fff?�u�?&찗d@T�����?�`?U?ȩ?X���� Z���T:z�TB��Wa� з*dů�ρϺϥ��� �����&�8�#�\�h�+�F. Kߘ�G߼��3���Wɯ���G�@ G����X� C�|�g�y������� ��jZ���ￏQ��� ��ߙ�����3����� ��/A��t_P�������� ���b���@+�Fp�IP�t��2%���[`B�0����<ze�cb!�@I�
�M`B�@��@`�9�@y��?�h�� �@�3��[N��N�N�E��<�/:/�L �>��ڟ��A�p�C�F�@�S�b/DpX������@�t��%�h��`/�qG��Gk�nF&�Fצ�pE,8{�/ �F�ZG����F�nE�D�E,ڏ�/� ����G��F7���F��ED�� .��C?.?g?R?d?�? �?�?�?�?�?	O�?O ?O*OcONO�OrO�O�O �O�O�O_�O)__M_ 8_q_\_�_�_�_�_�_ �_�_o�_7o"o4omo Xo�o|o�o�o�o�o�o �o3WB{f �������� �A�,�Q�w�b����� �����Ώ���=��(�a�L���p�����(�r!3�ji��r��y�ꕢ�3Ա�ڟ<�y�4 ����y��P�2�D�&��jb^�p�1w���������ʯ@���ܯ� �s�P^�	PD�c�`�m���y� \������Ӱ�¿Կ �����.�G�� ��}ϳϡ���홍�U� _�J���$�y.�@� v�d�z߈ߚ�x�4�ހ������ ��D�.�2v� �$[�G�[Ϣ^�B���B��CH� ^����u���� �������p�h�M�@_�q����������E^�^�Y�m�2��
 ����# 5GYk}�������h*�� ���>�x}��$M�SKCFMAP � ���� ����m�N"ONREL  6��9_�"EXC/FENBk
7]΄FNC�}JO�GOVLIMkdtuyd"KEYku�"RUN���"SFSP�DTYU��v_S�IGNk}T1M�OT�z"_C�E_GRP 1n��9\���/�� �/�/4��/?�/2?�/ '?h??�?C?�?�?y? �?�?�?O�?@ORO	O vO-OoO�OcO�O�O�O _�O*_<_#_`_-�"�TCOM_CFG 1o/���_�_��_
|Q_ARC_�6��UAP_�CPL�_�NOCHECK ?/ 5�;h9oKo ]ooo�o�o�o�o�o�o��o�o#5GTN�O_WAIT_L�F'5y"NT�Qp�/���q_ERR�!2q/_��  R_���"�:��L�dT_MO�sr>�}, 7�P_���_�PARAM�rs/������MW��� =e�345?678901.�@� R�)�q���_�����˟`����ݛLW�3��E�؏i�cUM_RSPACE,��������$ODRDS�P�SI&�OFFSET_CARTo�ݨDIS�ݢPE?N_FILE�I!��Q�v�POPTIO�N_IO���PW�ORK t�'F� T�|�
� ^�F� �
���Z���	 �m���A�
���i�_DSBL  ��v���ޡRIENTTOj�C���8�ῠ�UT_SIM_D�J�6	��VàLCT u�}\���Q��W�_PEXE���RAT����� ���UP ve����������Ϭ*�8��$��2�#h�)deX)dh�>O�X dY�� �ߣߵ���������� !�3�E�W�i�{��� ����������2n�� )�;�M�_�q���������<����� +=Oas����X��� O��1m(?���(�.�g�}�"0 �д�u�  @D�  &�?��?р~H�D4  Ez�Z3;�	l	� 0ӀS@(SM� �i�i ��H)!H,��H8�Hm��G�	{G�8��6�MV��� �SC�)���)�����Ճ�*  �_p  � > �� ,�//)/ �B,�Btr�«{�H�¼�/���/�"�# �,�0 �� �  �� ߽pj  B ��&X�?MU	'� � 12�I� �  ����-=���8U?g;/�@}?�0 ~.ѱ�?;Ѳ���rH[N5��?  'M�XD�> C)�f)�J BN +��=%O7O�R��@D1�o�o$����JWAD0�J5�4�: �1�E &?�O�O#__G_2]��� �t �O� ru �4 ��R<�Uɳ� :�%Ё�р� �?�fAf��@[�_�_V_{��o~��18р"o0j>�P�Q6YPрZo�W�rAdS�%�>L�w0�#�<	�I<�g�<#�
<�2��<D��<��׍�l�_��ѳMb�@?fff�?�0?&p:T@T��q?�`?Uȩ?X�-q �iyBq5Ya ��gI�_���� ��!��E�W�B�{� ��d�����ՏLnp�Ώ/�ʈG�@ G��U�ȏy�d����� ��ӟ�������yB =� ��?p���/򏸯 �߯R���'�9��o N�`�����~�����ۿ
ƿ�B�ĮD�e��ֿ;�ҿ_�J�?�A�h�oϨϓϸ��D4	��b!�_@���� �ħ��Ŀ����%�@I��)�M`B@���@`�9@y���?�h	� ��@�3�[N���N�N�E���<�/Y�kЖ�>��ڟ�A��p�C�F@��S���pX������@�t���%�h��߉!G���GknF�&�FצpE�,8{�� F���ZG���F��nE�DE,�ڏ��ૐ�G���F7��F?��ED��Mf�� b�M��q������ �����(��8�^�I� ��m������������� ��$H3lW� {������ 2VAS�w� �����/.// R/=/v/a/�/�/�/�/ �/�/�/??<?'?`? K?p?�?�?�?�?�?�? O�?&OO#O\OGO�O�kO�O�O�O�N(]�3g�ji�O�a��	U�E3Ա��O_<q�4 ��%_7_<q��P�Q_c_ERj�b}_�_1w������]�Y�_�_oP�_1ol��P�bPcn~���o�O�o{_�o�oY�`��o�o, /;M#�f0o�� ���Y�et�~�i#�1�C�yM�_����� ������{bS�Ԏ���	�?�-�c�Mj2����$�VG�z}�Bh����B��CH� }�9�֟�����0�B���wl�~��������Ư�T����\��qQ��U
 ί�0�B�T�f�x� ��������ҿ����܇��� ��]{x}���$PARA�M_MENU ?�Յ� � DEF�PULSE�	�WAITTMOU�Tl�RCV� �SHELL_�WRK.$CUR�_STYLj�Ϋ�OPT����PT�B����C��R_DECSNw�Te'�!� 3�E�n�i�{ߍ߶߱� ����������F�A��USE_PROG %P�%B��V�CCR��UeXÚ��_HOST !FP�!�����Tt`���������4���_TIME�� �T��  A�GDEB�UG��P�V�GINP_FLMSK]���TR����PGAʹ� |�[���CH�����TYPEM�Y�A�;�Qzu� �����
 )RM_q��� ����/*/%/7/ I/r/m//�/�/�/�/��/?��WORD �?	��	RS���CPNS�E̺�>2JO���BT�E���TRACEgCTL�PՅZ�� {`� �a`{`�>q6DT� QxՅ�0�0�D��Sc�{a�0���2��Q�?�?�2�4D1�2#A�O.O�@ORFcA�bB`D	�`D
`D`D`D�`D`D`D`D
`D`DObOtO�F A�5P�2Q0TOB�PRPBP�BP 0T�BP�BP�BP�A,_>Z�_=_O_a_s^ $_�_�_
b��"o4d�_ �_�_�O�O__a�1�	ad�TVd�^dfdnb�Wr�k}�o�o�j;qwc�TvT~T5Oc M_q�����v ,>�
�t�@�R� d�v���������+� �����ˏ��,�>�P� ̟ޟ���9�*� <�N�`�r��������� ̯ޯ���&�8�J� \�n���������ȿڿ ����"�4�F�X�j� |ώϠϲ��������� ��0�B�T�f�xߊ� �߮����������� ,�>�P�b�t���� ����������(�:� L�^�p����������� ���� $6�F l~������ � 2DVhz �������
/ /./@/R/d/v/�/�/ �/�/�/�/�/??*? <?N?`?r?�?�?�?�? �?�?�?OO&O8OJO \OnO�O�O�O�O�O�O �O�O_"_4_F_X_j_ |_�_�_�_�_�_�_�_ oo0oBoTofoxoN �o�o�o�o�o�o ,>Pbt��� ������(�:� L�^�p���������ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v����� ����п�����*� <�N�`�rτϖϨϺ�����$PGTRA�CELEN  ���  ��������_UP y���љ������_�CFG z�)������<���� <�Z�l�<�$�D�EFSPD {�/��a�����I�N'�TRL |�/�S�8Lԃ�IPE�_CONFI+�}>���<�]x�LID(�~/���GRP 1���������@��
=�[���A�?C�C
�XC)��B��r������dL�z�������� 	 �r�N��Ҩ�� ´����B������������A���> �6>7�D_�������� ='�=)���������	 B-��Q�M���  Dz����
��&L7p [�������/�6/!/Z/��
�V7.10bet�a1<�� B�=q�"`ff@���">����!=���͏!A>ff޷!@�ff�"�\�)�"D��?� � �!@�!� �!Ap�#W��h/??*?<?FK;�w����O/ �?K/�?�?�?�?O�? O>O)ObOMO�OqO�O �O�O�O�O_�O(__ L_7_p_[_m_�_�_�_ ��_ o�_$oo!oZo Eo~oio�o�o�o�o�o �o�o DQy{/�#F@ {yw}�y{ ջy�-������ /�Z?l?~?w���t��� ��я��������� O�:�s�^��������� ߟ�ܟ� �9�$�]� H���l�~����_ۯ� �����5� �2�k�V� ��z�����׿¿��� ��1�\n�j�|϶ �������	�4�F� X�j�c�χߙ߄߽� ���������)��&� _�J��n������ �����%��I�4�m� X�����ί�������� ��!E0B{f ������ H�Zό�Vh�ϴϊ ����� �2�D�V� O/�s/^/�/�/�/�/ �/�/�/? ?9?$?6? o?Z?�?~?�?�?�?�? �?O�?5O OYODO}O �O���O�OtO�O�O_ �O1__U_@_R_�_v_ �_�_�_�_�_"4F xBo|����o� �o�o//0/B/;�_ _J�n���� ���%��I�4�F� �j�����Ǐ���֏ �!��E�0�i��O^� ��N�ß՟������ �A�,�e�P�b����� �����o o2oTo.� hozo�o�����o��Ϳ �o
گ'�֯K�6� o�Zϓ�~Ϸ��ϴ��� �����5� �Y�D�V� ��z߳ߞ��������� �1��Uy��:� ���������	���-� �Q�<�u�`�r����� ������T�f� x�n�������� ����7"[F j������ �!//E/0/i/T/f/ �/�/�/�/�/�/?�/ /?A?l�e?w?&?�?�? �?�?�?�?�?OO=O (OaOLO�OpO�O�O�� ��*�O_@RdZ_�l_��$PLID�_KNOW_M � ����A�TSV �v��P�[?�_�_o�O&oo�#o\o�B��SM_G�RP 1��Z� d�I`�oo�$Cf�d����D��TPbj�oLk �f�o"~�U�o> n2T�~��� ��7�4���p�D� ��R���ʏ�������� ��6�
�T��*�����V�QMR�c��mT�EGQK? GR��(� #���[��/�A�S��� ���������$���� W��+�=�O������� ����� ���S�����ST�a1 1�j�����P0� @����E�ϲ��� ������M�0�B�T� fߧߊߜ���������@��7��,�m��2��9���A�<��z�A3�������4���������5)�;�M�_���6x���������A7����������8�(:L��MAD � ���� ��P�ARNUM  ��Ko���SCH
�
 �
��S+UPD��xaq|{��_CMP_�`�� <Pz '�U�E�R_CHK��a��Z���RS���_�Q_MO� �%�_��_RES_G����� ��v/ {/�/�/�/�/�/�/�/ *??N?A?r?e?w?J'��W,g/�?L%��? �?�?N#(��?OON# w�4OSOXON#��sO�O �ON# �O�O�ON#d ��O__N"V 1�x�Uua�@cX��P}p�P$@cW،P}��P@@cV��P��"THR_IN�R���pbA%d�VM�ASS�_ Z�WM�N�_�SMON_QUEUE ��eT��`Ȩ`�N��U�N�V�2`ENqD4a6/NiEXE]o�NeWBE\`>o/cO�PTIO;g?+2`P�ROGRAM %j%1`O_�0b?TASK_I��nOCFG �ox�9pDATAɓ]�B{@ev2w� �����z��+� =�O��s���������^nzINFOɓ��}�!dr��!�3�E�W� i�{�������ß՟� ����/�A�S�e�w�4҇ބ��| �98q~�DIT �B|ׯj~WERFL~h�wS~�RGADJ {�ƪA�  ,��?E�8��Q�IOR�ITY�W���M�PDSP�a�j�U��WvT�OG��_�TG���Rj��TO�E�P1�ƫ (/!AF�PE5 �~��!tcp��>%�!ud�?�!icm<�Q_���XY_<q�Ƭ=�Oq)� *������Op��������� ���<�#�5�r�Yߖ� }ߺ��߳������&�=*�PORT�a��OpA%�_C?ARTREP~`Ʈ>��SKSTA�X!*�SSAV`�ƪ	�2500H80A9u�T毙䕣�ƫ�����`X#�x$�6�m�URGEU`�B��A)WFP�DO�V�2�W�q�?Q��WRUP_DEL�AY �Ưe�RO_HOT�hwR%z�����R_NORM�AL�n��6SE�MI:y�QS�KIP���X%�x 	����� ���X%-;% [mE���� ���!//E/W/i/ //y/�/�/�/�/�/�/ ?�/?A?S?e?+?�? w?�?�?�?�?�?O�?�+O=OOO1U�$RB�TIF��NaRCV�TM�����m@DkCR����A�@�u�B��r�A�U���@�-߃)�����{�;/ž؞~�Ꮹ�_��_ �<	�I<g��<#�
<2���<D��<��
+__{_�_)`���_ �_�_�_�_ oo$o6o HoZolo~oi_�o�o�o �o�o�o�o DV �_z������ �
��.�@�R�=v� a�����������׏ �*�mN�`�r����� ����̟ޟ����� 8�J�5�n�Y���}��� ȯ�����A�"�4�F� X�j�|�������Ŀֿ �ӯ���0�B�-�f� Qϊ�m��������� ��,�>�P�b�t߆� �ߪ߼ߧ�������� (�:�%�^�A����� �������� ��$�6� H�Z�l�~���{���� �������� 2V h������� �
.@R=O �s�����/ �*/</`/r/�/�/ �/�/�/�/�/??&?�28�AGN_ATC� 1��K �AT&FV0E�02;ATDP�/6/9/2/9�p8ATA2>,�AT%G1%�B960k9+�++�?,�1H�?,��AIO_TYPE'  EC/4?�REFPOS1 �1� K x�O[H/O/�O�M NO`O�O�O�O_�OC_��Og__d_�_+K2 1� KLON_�_o��_*o�_5A3 1� �_�_�_ o�o�o�o@oS4 1�Woio{o�o3W�oS5 1��o�oJ��|�jS6 1������]�H����S7 1��(�:�t���ݏ���S8 1�����Ϗ	���r����)�SMASK 1� O  
���ɗ'XNO�?���1.��8�1AMOTE  ��.DN�_CFG ��U���5�0BPL_RANGQ�K!Y��POWER ��Q5 a�SM_D�RYPRG %��%R���ȥTAR�T ����UME_PROׯ�d��.D_EXEC_E�NB  �5]�GSPD=����Y3��gTDB����RMÿ.��MT_ѐT��S��D0OBOT_N�AME ��S�;9OB_ORD_NUM ?���AH80�0I$�	��se	�\������ ��e��	@��}�D|��D0PC_TIMEOUT��{ xD0S232n��1�Q; L�TEACH PE�NDAN��j�5���=Q�x0Mai�ntenance ConsK"-���"+�t4KCL/)C�}�6��|�� No Us�e�=[߹�F���NPqO�ќ�5�_����CH_L@���U���	J��MAVAIL`���+���]�I�SPACE�1 2�=L �����p��扢�J@����8�? ��� ���V�w�N� �������������� 4�&G
l�}d	Q5 U1���������` 4&G
l}d�#��2������ ��2A/b/%/w/�//�/�3��� �	/�/-/O/^??B? �?�?�?�?�4�/�/ ??&?�?J?l?{O�O@_O�O�O�O�O�5�? OO1OCO�OgO�O�_��_|_�_�_�_o�6 _*_<_N_`_o�_�_ �o�o�o�o�o!�75oGoYoko}o+�o �o����)��>��8Rdv��H� ����ӏ%�F�-��[��G ��� R�;�
�� ����ԟ���
�� .�@����c���p���8�¯=�dؠ��ϟ�� �!�3�E�W�i�_�q� �����x��կ�� '�9�K�]�oρ�w��� ����Ͽѿ����5� G�Y�k�}ߏߡߗ���p������� `S� @��8堯F�"�*ل������ �������,���� V�h�2�<�N������� ������.L4 v�R\n�����
f�7�_MO�DE  ��MS ���&����AÏb��*	��&/�$CWORK_{AD]	3��!/R  ���t �+/^ _INTVA�L]���hR_O�PTION�& �h�$SCAN�_TIM\.�h��!R �(�3�0(�L8������!��3��1��/@>.?����S22�41�9dD�4�1"3��@��@�?�?�?���IP���@���JO8\OnOE@D���O �O�O�O�O�O__(_�:_L_O���4�X_�_�_��8�1���;�o�� 1��p�c]�t��D�i�1��  � lS2��15 17oIo [omoo�o�o�o�o�o �o�o!3EWi {����wc�� �	��-�?�Q�c�u� ��������Ϗ��� �)�;�M�_���`[ ����ğ֟����� 0�B�T�f�x������� ��ү�����$�7�  0��� om�� ������ǿٿ���� !�3�E�W�i�{ύϟ� ��������v���/� A�S�e�w߉ߛ߭߿� ��������+�=�O� a�s�����ߖ��� �� ��$�6�H�Z�l� ~���������������� 2DVP�\�  �A������ �%7I[m �������/ �/C(/N/ `/r/�/�/�/�/�/�/�/?F;/?B?F;�x1 ;?w=�	123456�78{��
l�@�P�?�?�?�?�?O9/2ODOVO hOzO�O�O�O�O�O�O -/
__._@_R_d_v_ �_�_�_�_�_�O�_o o*o<oNo`oro�o�o �o�o�_�o�o& 8J\n���o� �����"�4�F� X�j�|������ď֏ �����0�B�T�f� ����������ҟ��� ��,�>�m�b�t��� ������ί����(��6yI�[�@�`����������Cz � Bp*   ���254F��$S�CR_GRP 1��(�e@(�l߀�0@� `1 �[1s	 )�3�C�<�t� vrY�8P�}�kϤ�n���95C�����-u��ȡ����LR Mate 200iC �1�90�1Շ0LR2C �3�=OÆ�ED�
f؜1u�2�@U7��`1��v��@�u���	t��������4�$�^0�2��� _2T�gϡϊ��o�F� D�f?��s�����￶}ht ,Z�qO� -LN�B�˰�P�N��g�N�Aܰv�  @�DЎ�N�@����  ?� ��J�H˰��y��N�F@ F�` ������A,Q wb���n�N���������B� �_J�n�� ���/�%//I/ ��E+:3��6?|?�5�ա
�/�/�#��@=���"�/pǢ� 3Bm�07�590@7����EL_DEFAULT  I���� �^1MIPOWERFL  V�v5]2΃0WFDE�m4 �v5 �ERVENT? 1���O�t3�C�L!DUM�_EIP?�8�j�!AF_INExj0O�$!FT�?�=NOaO!Q�O ��PO�O!RP?C_MAIN�O�Hq��O�O�CVIS�O�I��OE_!TP&8PPU<_�9d4_�_�!
PMON_POROXY�_�6e�_��_XR�_�=f�_)o!�RDM_SRV�*o�9gouo!R�R8�o�4hdo�o!
��@M�_�<i�o!RLSYNC�4y8�oY!R3OS�?�|�4H� tO�8c����� ;��_�&���J���n� �����ȏڏ7�I���m�4���X����7I�CE_KL ?%��; (%SVCPRG1���안�!��3*�/��4�R�W��5z���6�����7ʯϯ�C�$�5�9��o G����o������ D����l��񑔯� 񑼯7���_��� ���4����]���� �������'��տO� ���w��%ϟ��M� ���u�������� ��?�A��Ͽ�ђ�؟ ꐊ���ɱ������� �?�*�c�N������� ����������) ;_J�n��� ���%I4 mX�|���� �/�3//W/i/T/ �/x/�/�/�/�/�/�/�?/??S?Ś_DE�V �9��MC:[8�i.m4OUT_Rf1~6~i8REC 1����f0�0 �1 	 �2�?�1���3O�MO@O+OdO��
 ��Z���6 �s  UEBf0KX�q�0�0�f0ʬ��2�3f0nf0�@ ���-�X�O�2E0��0'qE0_�O_�5 "_�C&_L_:_p_^_�_ �_�_�_�_�_�_o o "oHo6oloNo`o�o�o �o�o�o�o D 2TVh���� ����
�@�.�P� v�X�������Џ��� ��*��N�<�r�`� ������̟��ܟޟ� &��J�8�n���b��� ��ȯ��دگ�"��3 ~A�(��P���t��� ��ο�¿��(�� 8�:�Lς�dϒϸϦ� ���� ���$�6��Z� H�~�lߎߴߢ��ߺ� �����2� �V�D�z� ��n���������
� ��.�@�"�d�R���v� ������������ <*`N��x� ����8 HJ\�������G�5V 1��< �P_�1�GFO�2�  jH�0wXJ>a?_TYPE�?k2�HELL_CFG� �z:f2/ ��B�/�/ %RSR�/�/�/?
?C? .?g?R?�?v?�?�?�?��?�?	O�?-O?O/�  �!�@oO�OP�O�C�I�AP�OL�B�@�WgB2P�d�O�O�&HK 1��+ �OE_@_ R_d_�_�_�_�_�_�_ �_�_oo*o<oeo`o�ro�oa&�#OMM ���/�o�"FTOV_ENBr$!}*�OW_REG_U�I�oe"IMWAI�T�b�I${OUTrv$&yTIMuw��`VAL5>'s_UNIT�c�v�})MON_ALI�AS ?e�i ( he!� �� $�6�Q&�c�u����� D���Ϗ�����)� ;�M�_�q�������� ˟ݟ����%�7�� H�m������N�ǯٯ ������3�E�W�i� {�&�����ÿտ習� ��/�A��e�wω� �ϭ�X��������� ��=�O�a�s߅�0ߩ� �����ߊ����'�9� K���o�����b� �������#���G�Y� k�}���:��������� ��1CU y ����l��	 -�Qcu�2 ������/)/ ;/M/_/
/�/�/�/�/ �/v/�/??%?7?�/ [?m??�?<?�?�?�? �?�?�?!O3OEOWOiO O�O�O�O�O�O�O�O __/_�O@_e_w_�_ �_F_�_�_�_�_o�_ +o=oOoaosoo�o�o �o�o�o�o'9 �o]o���P�������s�$S�MON_DEFP�RO ����:� �*SYSTEM*  �l�*��RECALL ?�}:� ( �}�5xcopy f�r:\*.* v�irt:\tmp�back��=>l�aptop-u9�nqdgeh:5�928 ��3 723 5�͏ߏ�s}6z�a���������B�T��:{�s:o�rderfil.dat������ӟ��}1{�mdb: �������=�O�a�� y�������ү��� ����-�>�P�b�u��� �����ο����� )���L�^�q����� 9���������%����H�Z���
xyzrate 61 �@�)�;�������!z�~��39020 ����?�Q�c���tp?disc 0����,��������t�pconn 0 ������J�\���; z������6�������2������>Pb ��ߕ��1��g7�ϋ��DV i�{������g ����@/R/d/w 
/��/�/�/��/ �/+<?N?`?s�/ �;?�?�?�?�?'/ �?JO\Oo/�/?�/7O �O�O�/�/�O#?�OF_ X_k�}�_!_3_�_�_x�����7068���_=oOoaot�{B�So�utput\ca�lpr.pc�0:� over =>�33554432:100017��2o�o�ohN3zhtemp�joc�o?Q�c��4zotest.ls�o�g/��0�w5�p�rtp~� ��s�H�Z�m��f �,���Ϗ���� ���M�_�r?�?Ok 6�ǟٟ�?�?��h�� >�P�b�uO�_�(t2��ïկ�O�O����8  ��C�U�h�z����0� ��ӿ��������?��Q�c�  �$SN�PX_ASG 1߶������� P�'�%R[1]@g1.1f�l�?��s%���Ͽ� �����6� �@�l�Oߐ�s߅��� �������� ���V� 9�`��o������ �������@�#�5�v� Y������������� ��<`CU� y������& 	0\?�cu� ����/�/F/ )/P/|/_/�/�/�/�/ �/�/?�/0??%?f? I?p?�??�?�?�?�? �? O,OOPO3OEO�O iO�O�O�O�O�O�O_ �O _L_/_p_S_e_�_ �_�_�_�_ o�_�_6o o@oloOo�oso�o�o �o�o�o�o V 9`�o���� ����@�#�5�v� Y�������Џ��ŏ� ��<��`�C�U��� y���̟���ӟ�&� 	�0�\�?���c�u��� �����ϯ���F��)�P�|�_�x�PAR�AM ������ �	���P���p�OFT�_KB_CFG � ����״PIN_SIM  �ˁ̶�/�A�ϰx�R�VQSTP_DS�B�̲}Ϻ���S�R �	�� &� TEST V����ԶTOP�_ON_ERR � �����PT�N 	���A��RINGo_PRM�� ���VDT_GRP �1�����  	 з��b�t߆ߘߪ߼� �������+�(�:�L� ^�p��������� �� ��$�6�H�Z�l� ~���������������  2DV}z� ������
 C@Rdv��� ���	///*/</ N/`/r/�/�/�/�/�/ �/�/??&?8?J?\? n?�?�?�?�?�?�?�? �?O"O4O[OXOjO|O �O�O�O�O�O�O�O!_ _0_B_T_f_x_�_�_ �_�_�_�_�_oo,o >oPoboto�o�o�o�o �o�o�o(:L sp�������� ��9�6�׳VP�RG_COUNT������d�EN�B/�_�M��鴖�_�UPD 1�	�8  
M������ �-�(�:�L�u�p��� ������ʟܟ� �� $�M�H�Z�l������� ��ݯد���%� �2� D�m�h�z�������¿ Կ����
��E�@�R� dύψϚϬ������� ����*�<�e�`�r� �߭ߨߺ�������\�YSDEBUGn��Ӏ���d��"�SP�_PASSn�B�?4�LOG �V΅�������
�  �����
�MC:\`��a�_MPCf�΅����ҁ���� ҁ��SA/V �i��������SV�T�EM_TIME �1�΋ (u���q�������T1S�VGUNSɀo�'������ASK_?OPTIONn�΅�������BCCFG �΋O���I�2��`;A�I�r ]o������ �8J5nY� }�����/� 4//X/C/|/g/�/�/���,�/�/ ??�/ �/H?3?l?W?�?��? ��0�?�?�?O�?&O OJO8OZO\OnO�O�O �O�O�O�O_�O _F_ 4_j_X_�_|_�_�_�_ �_�_o�X�  o2oPo boto�_�o�o�o�o�o �o�o:(^L �p����� � �$��H�6�X�~�l� ����Ə���؏���� �D�2�h�o������ ԟR�����.�� R�d�v�D��������� �Я����<�*�`� N���r�������޿̿ ��&��J�8�Z�\� nϤϒ���~������ "�4߲�X�F�hߎ�|� �����ߤ������� B�0�R�T�f����� ����������>�,� b�P���t��������� ����(��@Rp ������� $6ZH~l ������� / /D/2/h/V/x/�/�/ �/�/�/�/
?�/?? .?d?R?�?>�?�?�? �?�?r?OO(ONO<O rO�O�OdO�O�O�O�O _�O__&_\_J_�_ n_�_�_�_�_�_�_�_ "ooFo4ojoXozo|o �o�o�o�o�? 0 BT�oxf��� ������>�,� b�P�r�t��������� Ώ��(��8�^�L� ��p�����ʟ��ڟܟ �$��H��o`�r��� ����2�دƯ�����2��P��$TBC�SG_GRP 2���� � �P� 
 ?�  {���w��� ��տ��ѿ���/�A��T�[��b�d0� �p�?P�	 H;BHA�L�͌�@�B   C���϶˘���ϟ�D����AQ���x���A��T$��9��6ff��f�@2P�C�ώ�@�f߬��C��ߐ߮ߴޥ� ��%��%�D�W�"�4��j�|�������?�Y�����	�V3.00s�	�lr2c��	*�2�*�O�A� ��ѳ3e3P�d��� x�J�y�  �������T�JCFG Ė�l� o������������=K
%�Kq\ ������� �7"[Fj� ������!// E/0/i/T/f/�/�/�/ �/�/�/s���??(? �/[?F?k?�?|?�?�? �?�?�?O!O3O�?WO BO{OfO�O�OP�<��O ��O�O�O0__T_B_ x_f_�_�_�_�_�_�_ �_oo>o,oNoPobo �o�o�o�o�o�o�o :(^L���� ��h� ��$�� H�6�l�Z�|�����Ə ��֏؏� ��D�V� h�z�4�������ҟ ԟ��
�@�.�d�R� ��v��������Я� ��*��:�<�N���r� ����̿���޿ �&� �>�P�b�ϒπϢ� �϶��������4�F� X�j�(ߎ�|߲ߠ��� ��������B�0�f� T��x�������� ���,��P�>�t�b� �������������� &(:p^�� ��t�����6 $ZH~l��� ����/2/ /V/ D/z/�/�/�/j/�/�/ �/�/?.??R?@?v? d?�?�?�?�?�?�?�? OO<O*O`ONOpO�O �O�O�O�O�O_�O_ _&_\_�t_�_�_B_ �_�_�_�_�_"ooFo 4ojo|o�o�o^o�o�o �o�o�o0B�o xf������ ���>�,�b�P��� t���������Ώ�� (��L�:�\���p��� ��ʟ��� ��_�*� �_�l�Z���~����� į�د� �2��� h�V���z���¿Կ� ��
�����.�d�R� ��vϬϚ��Ͼ���� ��*��N�<�r�`߂� �ߖ��ߺ������� 8�&�H�n�\���>� ����x������4�"� X�F�|�j��������� ������
Tf x�D����� �P>tb �������/ /:/(/^/L/n/p/�/ �/�/�/�/ ?�/$?6? ��N?`?r??�?�?�? �?�?�?�? OODOVO hOzO8O�O�O�O�O�O��N  PS �V$_R�$TB�JOP_GRP �2��E�?  ?�W<R�CS�J\��@�0WP�R@T�P ט ��T�T ��Q[R	 �BL�  �UCр D�*W[Q�_�_?ff�fe:lB ��P�ff@`�?33D  $a�U 3o>g�_�_po�l�P�e�9<�bbY���?٪``$o�oUAm��gD�`$�co�Quz9�P��Aa�P@a����C�Z`Ep�o]A63ffpu`aD/�U�h�͔r��~�a�R@ieAq�`�q��@9q�|�d&`%���c�333D�\P8���?�`?L�pAp[QB�b�k�}� ��z>�� >�ffԁL���T�f��fo � �Nw@�*�8�f���r� ,���П��ȟ��'�� ��F�`�J�X�����S�C�Vء��	�V3.00�Sl7r2c�T*��T�Q�� E����E�A E���E��3E��iNE�!hE��فEۑ�E��I�E��E����E�rF��F�F�M(F�5F�BFaOF��\F"f,�z�  E�@ E��� E�� E��  E����� �E����� E�ꆰԎ�ᆰ� �F   F� �F$ Fj` �F�@ F�P �F�` 9�IR/9�o���L�Q_ ��V���LQ�8TESTP�ARS�XUP9SH�Rk�ABLE 1%�J[4�SV�+�Q �0�V�V�VȨWQV�	V�
V��Vȥ�QV�V�8V�뱅�RDI��TQ�϶���������f�On߀ۊߜ߮�������Sl�RS 0ړ�� �����������#�5� G�Y�k�}��������� ����/]k�o��*	� %�7�I�����+�=��O؆�NUM  ��ETQ�P�P �밆�_CF�G ����Q@�<PIMEBF_T�Tq��RS~�;VE�R�<Q;R {1�J[
 8��RP� �@5  ������/ /&/8/J/\/n/�/�/ �/�/�/�/#?�/?Y?@4?F?\?j?|?{_��h@R
<PMI_�CHANG R >�3DBGLVQ`I�R;Q�0ETHE�RAD ?�E
;@�S �?�?TO6V��0ROUTe!�JZ!�D�OwLSN�MASK0HRSAA255.�E��O�O�8TOOLOFS_�DIq��5IOR�QCTRL �s[���n]8]_�_�_ �_�_�_�_�_o"o4o�Fo�
�_Tofo�og�PE_DETAIH�3ZPON_SVO�FF)_�cP_MOON �"P2�i�STRTCHK ��J^mO�bVT?COMPAT�h;C��d�`FPROG %JZ%j�=?~qqISPLAYr���j_INST_M��@ �|�g�tUS8e]orLCK��{QUICKME�0�)�orSCREF�}3Jtps��@or�a�f��2w�_{����ZyISR_GR�P 1�JY ؛ 6���@��;�)�_�M��8 ����Y�������͕ �����/��S�A�w� e�������ѯ��������=�+�M�s�	�12345678h����f�X`�1�Ћ�
 �}ipn�l/۰gen.htm�����0�B��X�Panel� setupF�}�<�ϘϪϼ����� u�k��*�<�N�`� r��ϖ�ߺ������� ��ߝ�J�\�n�� ����I�?������ "�4�F���j������ ��������_�q�0 BTfx��� ����>� bt����3�~�UALRM�pG {?J[
  � */!/R/E/v/i/�/ �/�/�/�/�/�/??�<?�SEV  ��n6�ECF�G ��m�6��A��1   Bȩt
 =?�s3E�?�?�? OO+O=OOOaOsO�Oh�Gz1ʂ��k S(Ο�OH7Isv?}{�`(%0?"_p_I_4_ m_X_�_|_�_�_�_�_��_o�_3o�L� ��M�OAoI_E�HI��p1��i  �(p ��(/�SOFTPART�/GENLINK�?current�=menupage,153,1}o0�o&�'�o�n71�oq���6qy);�eedit�b�T��`�	��-� �)oS�e�w������� <�я�����+��� O�a�s�������8�J� ߟ���'�9�ȟ]�@o���������è�R� �aR����%�7�I� L�m��������ǿV� ����!�3�E�Կ� {ύϟϱ�����d��� ��/�A�S���w߉� �߭߿���`�r��� +�=�O�a��߅��� ������ʯܯ�'�9� K�]�o�r�������� ����|�#5GY k}����� ��1CUgy ������	/ �-/?/Q/c/u/�// �/�/�/�/�/?��� ;?M?_?q?�?�?�/�? �?�?�?OO�?7OIO [OmOO�O�O2O�O�O �O�O_!_�OE_W_i_ {_�_�_._�_�_�_�_ oo/o�_Soeowo�o �o�o<o�o�o�o +?(?as��� ��o����'�9� ��o���������ɏ X�����#�5�G�֏ k�}�������şT�f� ����1�C�U��y� ��������ӯb���	���-�?�Q�<��$�UI_PANED�ATA 1������� � 	�}/f�rh/cgtp/�wholedev.stmc���ӿ�|���)pri��.�Ip}2�V�h�zό��ϰ� )���Ͻ��� ���0��T�;�xߊ� q߮ߕ��������Bv�Nq*�=�B� T�f�x�������3� ������,�>�P��� t�[������������ ��(L3p�i�� ������� ��1C�g �������L 	///?/&/c/u/\/ �/�/�/�/�/�/�/? �/;?M?���?�?�? �?�?�?0?Ot%O7O IO[OmOO�O�?�O�O �O�O�O_�O3__W_ i_P_�_t_�_�_�_�_ Z?l?o/oAoSoeowo �_�o�o O�o�o�o +�oO6s�l �������'� 9� �]�D����_o�o ɏۏ����#�v�G� �ok�}�������ş,� ������C�U�<� y�`�������ӯ���� ޯ�-�����c�u��� ��������T��� )�;�M�_�q�ؿ��|� �Ϡ����������7� I�0�m�Tߑߣߊ��� :�L����!�3�E�W� ��{�� ϱ������� ���r�/��S�e�L� ��p������������ =$a����}�r�����)�*��Vhz ������� �.//R/9/v/�/o/ �/�/�/�/�/?��������$UI_PA�NELINK 1����  ��  ���}1234567890_?q?�?�?�? �?�4��]?�?�?OO 1OCO�?gOyO�O�O�O��OYIY0:�M���[0-/SOFTPART/GENA1�?CONFIG=�SINGLE&P�RIM=mainedit �OI_[_�m_YJ_$_M=wi?ntpe,1@_�_�_�_XK  �_$o6o HoZolooo�o�o�o �o�o�o�o
2DV hz����� ���.�@�R�d�v� �� �����Џ���~�M 0,M9P� E=Por?S�,Ico:�{�^��� ����˟ݟ������7��[�m�P�������O���BS0ߢ��C���/�%�7�I�[�m� `C�������Ϳ߿� ���'�9�K�]�o��L ���э͙�Q|����� �����!ߨ�;�M�_� q߃ߕߧ�6������� ��%��I�[�m�� ���2���������� !�3���W�i�{����� ��@�������/ ��Sew���� .���z�!E (W{^���� ��/�//A/���� �Ϸ�}����/�/�/�/ �/?�2?D?V?h?z? �??�?�?�?�?�?
O O�ϝϯ�dOvO�O�O �O�OE�O�O__*_ <_N_�Or_�_�_�_�_ �_[_�_oo&o8oJo �_no�o�o�o�o�o�o io�o"4FX�o |�����e� ��0�B�T�f���� /���������ُ� ��>�P�3�t���i��� ��Ο��O/�s/(��/ L�^�p����������? ܯ� ��$�6�ůZ� l�~�������#O5OGO �� �2�D�V�h�� �Ϟϰ�������u�
� �.�@�R�d�v�ߚ� �߾������߃��*� <�N�`�r����� ���������&�8�J� \�n������������ ����m�"4ßXj M�q����� �BT7x� �����A��// ,/>/P/C�t/�/�/�/ �/�/�/o/??(?:? L?^?Ϳ߿�?�?�? �?�? OO�?6OHOZO lO~O�OO�O�O�O�O �O_�O2_D_V_h_z_ �_�_-_�_�_�_�_
o o�_@oRodovo�o�o )o�o�o�o�o* �oN`r��� ��m��&�8�� \�n�Q���u���ȏ�� ����"���?�?��{��$UI_PO�STYPE  ��5� 	�k�{��_QUI�CKMEN  �j�����REST�ORE 1ו5�  �A�/
�2�D�h�mc� ������¯ԯw���
� �.�@��d�v����� ��W���˿ݿO��*� <�N�`�τϖϨϺ� ���ρ���&�8�J� ��W�i�{��϶����� ���ߡ�"�4�F�X�j� ��������ߋ� ���y�+�T�f�x��� ��?����������� ,>Pbt��� ���(� L^p���I���� //��SCR�Eܐ?��u1sc-�u2�M$3M$4M$5M$6�M$7M$8M!��US#ER/ 4/F"T. O#SksW#�$4�$5�$�6�$7�$8�!��N�DO_CFG m؜�  ,� ��PDATE �)��None� V��SEUFR�AME  
���&,1RTOL_A�BRT7?��N3EN�BX?I8GRP 1��!��Cz  A��3�1��?�?�?�?�?FO"OG:ې�Ux81g;MSK � {5�Ag;N41�%a��B%��O��V�ISCAND_M;AXyEI�c8�@�FAIL_IMG�y@f���#�8�@IMREGNUMyG9
�KRSIZyC,����$,SONOTMOUW0{D�%��VU�#�c��� �P�2FR�:\�O � �MC:\XS\L�OG�VB@4 �!�O�_�Q�_o
�z MCV�_��SUD10fEXD9k
�f�wV�2ۜ���p(��=����o��j�o�o�o�o �o�o�o 2DV�hz��KPO64�_?S�0��n6�uQ0LI Q�z�x�q9V� �|f@�w��� =	�xSZV��~����wWAI���DSTAT 	ܛ;�@�_ď֏��$����EP12DW�P  ��P G/����q�AP-��B�_JMPERR �1ݜ�
  � 2�345678901�������ʟ��ϟ ��$��H�;�l�_��q����LT@MLOWp���P�@�P_TI_X��('�@MPHA�SE  53|��CSHIFTUB{1~k
 <�� �Ob��A�g���w��� ֿ���������T� +�=ϊ�a�s��ϗϩ� �������>��'�t��K�!��#ޛ:	VoSFT1�sV�@�M�� �5��4 ��0��UA�  BU8���Ќ�0p������Ҫ��e@��ME�*�{D�'���q��&+%�!�M�$�~k���9@�$~�TDI�NENDcXdHz�O x@[O��aZ��S���\�yE����G� ���2�����������RELE�y?w��^_pVz�_ACTI�V���H��0A ���K��B#&��RD��p��
1YBOX c��-�����2�D�19o0.0.� 83�;�254���2�p�&���robot��ԟ   �pN g�pc � �{�v�x�Ѽ�$%ZABC�3��=,{�낆;-!/ ^/E/W/i/{/�/�/�/ �/�/?�/6??/?l?!ZAT����