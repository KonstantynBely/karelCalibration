��   ��A��*SYST�EM*��V7.7�077 2/6�/2013 A�   ��	��BIN_CFG_�T   X 	�$ENTRIES�  $Q0FUP?NG1F1O�2F2OPz ?C�NETG  �D�NSS* 8 }7 ABLED? �$IFACE_�NUM? $DBG_LEVEL��OM_NAME �!� ETH_�FLTR.� �$�   ��FTP_CTR�L. @� LOsG_8	CMO>�$DNLD_F�ILTE� � SUBDIRCAP"n���HO��NT.� 4� H�ZA?DDRTYP� A =H� NGTHph���z +LSP� D $ROB�OTIG cPEEyR�� MASKa�MRU~OMGD�EVl%&�R�DM*�DIS���Y� TCPI��/ 3 $AR�PSIZoK_I{PFpW_MC-��F_IN0FA�~LASS�5H{O_� INFO���TEL� Pȟ���R WO�RD  $A�CCE� LV��$TIMEOUT�uORT �IoCEUS�  � ��$O#  �S���!��
��
� VIRTUAL�/��!'0 �%
U���F����04+5�'�� =���!�!j?����; x?�5��=2~;#"SHAR�� 19  Pf?O(4OHO7O lO/O�OSO�OwO�O�O �O_�O2_�OV__z_ =_�_a_s_�_�_�_�_ o�_@ooovo9o�o ]o�o�o�o�o�o <�o`#�G�k �����&��J� �n�1�C���g�ȏ�� 쏯��ӏ�F�	�j� -���Q���u����ן��ϟ0��7z _LI�ST 1�=x!1.k�09��j��1{��255.���r����05i�2 p���砖�����̯ަ3诂�_�� �2�D�ަ4`���װ��������ަ5ؿ��O����"�4�ަ6Pς���v�0�ϚϬ� �$��Q>�$% =� .6P+5U�o!R��)��0�H!� ����rj3_tpd���31 � �!!K�C� �߿�(�'6��!C� ;�����?!CON� ��z����smond���