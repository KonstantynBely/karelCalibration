��  ë�A��*SYST�EM*��V7.7�077 2/6�/2013 A�Q  �����ABSPOS_G�RP_T   � $PARA�M  �  �ALRM_�RECOV1   $ALMO�ENB��]ON�iI M_IF1� D $ENA�BLE k LA�ST_^  d�U�K}MAX�� $LDEBU�G@  
 ���APCOUPL�ED1 $[P�P_PROCES'0 � �1�����UREQ1 �� $SOFT�; T_ID�TO�TAL_EQ� �$,NO/PS�_SPI_IND�E��$DX�S�CREEN_NA�ME �SIGNj��&�PK_FI� �	$THKY�P�ANE7  	�$DUMMY12*� �3�4�G�RG_STR1� � $TIT^�$I��1&@�$�$�$5&U6&7&8&9'0''�%!'�%�5'1?'1I'1S'1�]'2h"GSBN_�CFG1  8� $CNV_J�NT_* �DAT�A_CMNT�!?$FLAGSL*�CHECK��A�T_CELLSE�TUP  P�� HOME_IO�� %:3MAC{ROF2REPRO8^�DRUNCD��i2SMp5H UTO�BACKU0 �� �	DEVI�C#TIh�$5DFD�ST�0�B 3$INTER�VAL�DISP�_UNIT��0_�DO�6ERR�9FgR_Fa�IN�GRES�!Y0Qy_�3t4C_WA�4��12HGX_D�#�	 d $CA�RD_EXIST��$FSSB_�TYPi� CHK�BD_SE�5AG�N G� $SLOT_NUMZ��APREV��|G �1_EDIT1_
 � h1G=�H0S?@f%$EyPY$OPc� �0LETE_�OKzBUS�P_CRyA$�4�FA^Z0LACIwY1�KR�@k �1COMM{ENy@$DGV�]QP� ���AL�*OU�B , C$�1V1AB0�~ OL�UR"2CAsM_;1 x�~f$ATTR���@0ANN�@�I�MG_HEIGH|yAcWIDTH��VTCYU�0F_�ASPECyA$�M@EXP;$ܸ Mf�CFcD ?X $GR� � �S!1U`BfPNFL�IC`~d
UIRE�s3��AOMqWI�TCH}cX`N.0S�_d�SG0 � 
$WARNM'@0f��@� LI? �a�NST� CORN���1FLTR�eT�RAT@0T�` ? $ACC�1"pp '|�'rORIkP�C�kRTq0_SF�� W �CHGI.1 [ Tz`u3IPpTYVD�@*
2 �P�`� 1zB*HD�SJ* ��qU2�v3�v4�v5�vU6�v7�v8�v9�u�qO�$ <� �so�o�h�s1�PO_�MOR. t� 0Ev�NG�8`TBA� 5c��@�A�����]@����ϋP�0Ѕ*��h�`
P�@�2� h�,p�J,p_Rr�rqo@+�J/r/�J�J	Vq@�Cj��m�g��lustP_}0OF� �2  @� RO_����WaIT8C��N'OM_�0�1ەq384 ��cD �;�d���hP���mEXp�G�0� F�p%r
�$TFx�JF�D3&ԐTO�3&@U=0��/ �H�24�KT1��E�� �e���f��f��0CP�DBG;a� k@�$�PPU�3�fc):��A�AX 1��dUN�$AI�3B�UFuF����! �|�`��`PI�U�Pr�Mq�M~��䠁�Fr�SIMQ�S��G��QE���"���MC{� �$�}1JB�`S�}1DE�C��������x� �ě0CHNS_E;MP�r$Gg�=��@_��q3
p1_FP󔞡TCh�@`�b���q0�c}�y�G�� V`�AԂ�!!���JR!0~ԂSEGFRA.p�v 7aR�T_LI9N�C��PVF������Y���Q���)B����( '���f�e�S���Q���.0�p�B��A����SCIZC�ћ�z�T���g������QRSINF3��p����?�������؉���Lot��G��*�CRC�eFCCC �`+���T�h��mh�Sb�A��h�*�f��:�DȬd�c��C��PTA�����w@�撀��EVT���jF��_��F��!N&�G�� X�������1i��! 1��,��hRGNP��"0qF���R}�D���2}�LEWN��Hc6����C�K�FA�dCx :�L��ou2��ԊA6N`Co�$L	Gp��B�1aP��s@��dWaA?@���~0R���dME%`��d��_RAs3dAZ�C���z�OkqFC�RH`X`F�`��}��,�ADI;�  6b� ���`�p�`5c�n�S�@1�7a�AMP$���PY8CU�Mwp�U��iQU� $ �P��C�CG1������DBPXWO��z��p$SK���2۱DBT TR%L�1 ��Q0Ti� �P�DJ�4LAY_CAL�1R !�'PL	3&@�0ED��Q5'�Q5'̡(�D�B��1!�W�PR� 
�1 0�1g" �PA$�q{$�� �L�)!#�/�#mp�0$�/�$�C�!%�/�$ENE�qr�&�/�#d R�Ep�"'H z�O)@"$LF3#$�#xB� W;���F�O[ _D0m�RO�(@���u��j���3R�IGGER�6PA�%S���ETURNܦ2RcMR_��TUr�`?�u0EWM���GN�P��zBL�A��E��$$P"#�CP� ��&@�Q"k�C5D�mpD�A#��p4\1i�FGO_A7WAY�2MO��fQ�g�CS_(<�QIS �����c�C���A�����B�t�Cn��A"�FW����DNTV@��BV kQ�����S˳W�sU��J&�U�� ��SAF�E�ZV_SV6bEOXCLUl�����'ONLA��SY��Q�tOTBa��HI_�V/M�PPLY_|�a��VRFY_#�q�Bd�_ )�0���_+�Ip ���@SG3� *�b݀�0 AM���a*����0��Vi.b%fANNUN� rLdKIDp�U�2~S@ �`mijarj�f`"p�OGI�"+��$1FOb�׀OT@w1� $DUMMAY���d[!�d١�|& �E, ` 8�HExs��b�SB�$�SUFFIA�@ ��@�a5�g�6�a�MSW�E-{ 8��KEYI����TMZ1^ӌq�1�v�IN����a!.{ D��HOST? !�r���t[ �t٠�tYp�pEM>���$�kR��pL��UL���/ �|3���;��DT50�!0 ϴ $9��ESAMP�ԕF���������I�0��$SUBe�Q�� �C�:��G�SAV��r����G�C� ˇ�PnfP$�80E��YN_Bn�1 0��DIadb�@O���}$]��R_I�� �E�NC2_ST � 2
ԇ J���L�q~S�`;����!3�M�I��1:�p�4  AL�3�M��0�0K�4x'a��AVER�q8��}�M�DSP�v��PC�U���\�ެ�VALUŗHE4� ��M�IP@����OPP7  �THS ���6�S�F�	F􁳠dL�0�T���SC�Q�d:�ET�o�5zrFULL_DUY�da�0��O�w�h�OT��A�0�NOAUTO�!6��p$�\���cTl�
�C!��C����۱�L�� _7H *�L���n�b���$�0P�˴ ��ֲ��[!���a��Yq���dq��7��8��9R��0����1��1��U1��1Ⱥ1պ1�U1�1��2
�2�����2��2��2Ⱥ2�պ2�2�2��3J
�3��3����3��U3Ⱥ3պ3�3��3��4
��-�v��SE�"8 <��~��`�;I�����/��FE�0�0� �9 ,��Q? z@^ ?�А��ER@#�q�A��z� :�`$TP��$VARI�B�:>��UP2�P; �pq�TD��S|��1`3���<�_B;AC�< T�pr���)��bP�P o�IFI)�P ���U���P��F�0��� =t ;'�Ԡ��P'�ST(&�� HR&�Pr0E����	%�C��	���_Cr�N�r��B���p�h�FORCE�UP%bn�FLUS
�`HN �E�h�R/D_CMK@E(����IN_��&vPg�REMM�F~Q���M �� 3
K	N0�EFF��N@sIN�A��OVMl	�OVAl	TROV̙��DT��mDTMX���m{@�
���? �*[ ��CL���_:p']@$�-	_�
�;_T��X
�J�@AQD� ��}���}!V1� RQ~��LIMIT_�ad椀�M��CLmd�}�RIV	�a��E�AR��IO*PC�C�����B�Bg�CM�@��R �GC3LF�G!DYM(/l�aR#5TWDG���| s%Ǵ�FSS& �s> P�a�!r1���wP_�!�(�!1R��E�3�!3�+5�&O�GRA���?w�i�kPW��ONT��EBUG)S&2*��P{@a�_E @� �p�P����TERMB5AK9O�RIG0BK5�0�GSM_�Pr�G0CK5�3�PTA�9DK5����UPB�Eg� -zAa�@.P|Y3.@A$SEG�:vf ELEUUSE�@NFI,��2�1xޠp4�4B$UF6P�$�FQ4@�wAG0TQ�&�HSwNST PATm�<piBPTHJ�AߠE�p��2�P؀	E)��؁��1R�@�InaS�HFT_��1oA�H_�SHOR ܣ�6 ��0$�7�@Dq�'�O#VR#�na�@I�@��U�b �QAYLO=�z��I'"�oAj�!�j�ERV��:Qh� �J��OG @�B0����U�>���R!P"�AScYM.�"��1WJG�уES�A�YvR�U�T @���E)�ᥳEaP!�WP!�WOR @�MB�� SMT�F�GR��3la�PA.@��jp�q�uG� � ����T�OC�1�`P�@ �$OP��ဝpՓá� ��O��RE�`RC�AO�pтpBe�`RmE u�h�A���e$PWR�IM�ekRR_�c�q�b.B H2H���p�_ADDR��H_LENGqByqnq�q��R��S�I H��S���q0Ӧu>Ӵu���u��SE�'�LryS��J $J�<�`��_OFF��r�PRM� �;�HTTP_�H��K (^pOBJ�?"ip��$��LE�`C!�ȠL � ��׬�AB_~T�S�s�S{`��*�LV�N�KR��eHIT���BG��LO�q t�fN�͂���`���`3SS{ ��HW��A��M�p`INC�PU�"VISIO �����+��t,��t,�~�� �IOLN���N̠�C��$�SLQb��PUTM_�$�`{�P x�V���F_AS�"O��$L��I���D�A��U�0�@Af��`q�<PHY���Ó�<���UO��#P `������ڔ� �2�pP���`(�L���Y�B�;�UJ�Q��z�NEWJOG�-G��DISx�<�K�-�f�#R 
�WAV��ǢCTR�CǢFgLAG�"[�LG�d�S ���Y�3LG_SIZo����������FD)�I �4�E�*��D0�� �c$���𖶦���K��D0��� SCH_ ��߅p�2��N��F�T���E�"~���D����U
�
�{`L�n	�DAU/�EA�0-��dE�;�GH�b;�BOO��Uh3 Aɒ��IT��y��[0ŖREC��SC�R��ʑDIēS.@��RGO���˒� ���d�´���SU����W�Ĳ�Ľ�JGM�$�MNCH,�F�NKEY%�KM�PRGK�UFY�PYطFWDY�HL��STPY�VY�@Y؀�Y�RS��H1`uۺ�CT���R��� �$�U	�m���
R�ݠғ2`�G=��@POd����Ŧ�M�FOCU�d�RGEX��TU%IK�I{�����	�@�����I�M��@A��S�`���@������A�NA���2�VAI�Ll�CL!�UDCS_HI+4`�s_�Oe�
!h�S���|�9S����IGN4���F�J��T�be�_B�Uj � V !PT�$*��rv�ϤT���AVrW !P�i�'���0�1?2�?3?d�__� X � i�=a�5��L�Ņ�ID� tbP5R��bOh ��\A�ST�	�RF�Y� �@�  _W$E�C�y����_�� Y L�؟0��@ ���`qFtǀ�Ft��Ѭ�_ Z ��p����b���>0C���[ �p CLD�P	��UTRQLI�{��T����FLG �� 1�O�D������LD���ORG������hW>(�spiT�r� 4\ �#0P��վ�Sy`T��70y ' �$�!�#RCLMC�$B/T/�)�Q��!=1I�p_d] �d�RQ73$DgSTB�p�   6l��-8AX�R /8�I<EXCES�b��`2Mp�1^�p@2�T�2��0_�p"6_A:&��;G?tY80K�d` \��GROU��t$M�B �LI9�CRE�QUIRDB�aLO�#KDEBUr� 1L
YM��agbʑ`@�4C�" 1ND��`�c`b���̨�CDC���IN'��C��Z`���H��N��a#�� �u1�APST�� �c\rLOC�R!ITp��P�Ap��1 1ODAQ��d� X�ON�cF �R�fV�	X��b�U����w �FX0I�GG�� e ��y X�a��X�XR�Q%��Y	��X	�x�V�0ғDATA�$`E�a�AS IN���f t $MDEaI:�)Sf��^d�![gH5P�@]ez��a_cANSW�a^d�a��^eD�)ARz�� nXpg �0CU4�qV�`�=URR2{�Gh D2�`A��A�!� d$CALI�&0��GS�w2K�R�INb�t<�INTEg�(i�bCu��X=RBqg�_N�qjPu�kr���$ht�2kuyDIV�&DHi0jp+�l $Vp�C�;$M�$Z0R<!�T 0R���b�em�H �$BELT|˪ZACCEL��q�;�"�IRCO��݁m��T���$SPSi0�Lt�ڰ�W��Cp8��T�9�P�ATH���.���3]��Pl1_<�r��Ł�"S Cr��_MG��$DD�9���$FW�`7`����.���DE�PP�ABNe�ROTS�PEEՂ@L� J�N�@��(0�t�$OUSE_p�P&�FܦSY>��p�! �Q�YN0A����OF�Fua��MOU߁N�GJ�܀OL~�ٔINC�d2Q��-2��<� -2ENCSpa`2U��+4R�IN��I]�B����"n�VE���s^�23_UP�օp�LOWL�� [�` '���D>�2 @Ep]'��2C[pW�gMOS���4MO���0�'PERCH  ��OV����蓼 ������$�8S+�� 2@������V�0^��O�L�P��7O�U�U�P"�������TRK|��AYLOA� J��1��]�͵³3P� ��RTI�1	�� MO�O�-2�28 �`4��wٳ��?�pD�UM2��S_BC?KLSH_C]�P� ϐΦ����bn�"�y�xÑ��!CLAL �V��!��� ��CHKt �SՐRTY�� ��C�
*!6a_�ä'_UM����C����SCL�W�LMT�_J1_L< 0-օa:�E4�U�G�D�8J�P�J�SPCd�ȑ�Z���3�PC �3�H�_A@���C� cX�T���CN_rN����.�S��%�V ���:����]�9���C' �SH�r� *�*!9�9� p��^����9���PA���_P��_�"�Ŷ�!ճ����JG����~��OG��,�TORQU��ON��޹*�B0٢-�*�L�_Wž��_�sj��sj��sj�I*r�I��I�sFKP]�aJ�!��c!�VC�0'42��1��{0��82��JRK��+~� DBL_SM��:�"M�@_DL�q�"GRVq�j�sj�s�KH_��I���
CcOS��LN-  �����p�	�p�	�����FZ� ٦KcMY�D�TH��eTHET0��N�K23�s��s� C-B�CB�sC&1n2������s��SB8�s��GTS�1W�C.�2Q�����$�<'3$DU���8�A!r�2P&�1Q�b8V$NE�4�PI � ���"%�v$�p��A��%�'���LCPH�5�"h��"S�� 3�33�"+3:2�pV�(V�(�p�,UV�*V;V;V";UV0;V>;VL9H�(@�&�2�-n�H;H;UH";H0;H>;HL9�O�,O�(O}I�.O��*O;O;O";O*0;O>;O2F�"��Y�T�'SPBA?LANCE_T@S�LE�H_�SP�Hq�hR�hR3PFULClX�R{W�R3�Uz1i
�UTO_<����T1T2�Y�2N���`��Tq����Ps d���T�O��p!�L�INSEG���REVf��Q�gDIF��zy1j_g6�r1k]�OBUa���t$yMI`���SL�CHWAR>��A�B��u$MEC�H�Tˑ�a��AX�˱Py��f�'�r�Pl� 
�bI��:�RO�B�CRW�-u�Ҷ-�MSK_KP��tn P �P_���R��r_tn���1 8�c�a�_p`�y�_p�a�IN:a�MTC�OM_C���po � ݀g`4�$ONORES��r��`޵rp 8U�GRlJ��eSD� ABג�$XYZ_DAx�!F�r�DEBU:aX�q���pq _P$��wCOD�� 1�����`��$BU�FINDXa� � !�MORRsr $�qU&���u��DӑyãHp"��bGi��s � $SIMUL��8��>����F�OBJEjP��A�DJUSψAY_I��8�D���s�nԐ_FIב=s�TZ��c����`b�"�(�b`p0G�D��F�RIW�d�Tg�RO�%�A�Eb�^�O�PWO> Vpt0>>�SYSBU0[�$SOP��I�����yU��b`PRUN�rڕPArpDٖ�b��.1�_OUTΑ�a��t$�IMAGҊ�\pv PDaIM���1�IN[ �0�RGOVRDY�˒����P�/�a�� L_`�PB�}����RB�ʇ ��MkᜪEDTb��` �N�@M��f~���]�SLjP�Vpu x $OwVSLfSDI��DEX���q�����$o��Vb��N�A�@�'��,�'�D�M~y��\�_SETK�Vpv @U�^��ep�SRI��j�
q�_��}�������dà*� �w H\q�`��A�TUS<�$TR�Cx T�X�ѳBTMTڷıI��P�4}Ѹ����Vpx D\pE���β�0Ehbϱ�8����ϱEXEհ�� ��)�=��f�ym�]pf԰UP�L�$�`6�XNN����������� �PG�uzWUBñ�e��ñ~��JMPWAI[��P���LO7о�F�A`��$RCVFAIL_Cwq����R9��p�c��(�}�"��-�AR_PL��D�BTB��,⾐BW�D ��pUM*�"�I�G�7��Qc�TNL�W�"�}�Ry�iӻ�E������Hp��DEF�SP` { L�\p�`��_��Ճ��UCNI����Ѐ�RD���Rb _LA`Pͱ��P�pUq|-�#��q��O��XPc�N�PKSET�
��Pq��Uq} h�ARSIZE5p��=��u��S̀OR��FORgMAT�Pg�COנ,q�<bEM�d�����UX��,��LI�b�Uq~  $>�pP_SWI�`V��/ G�b�AL_ )o���A�rB���uC�rD��$EL����C_lі� ?� � ���r���J30 �r��TI�A4Z�5Z�6�rMOM��f��s����pB��ADf��s�l����PU�NR����s�����ѡ��Rt�� A$PI�& E�kqE�p-~-� -�WC�0$��&¹�9q�gE��eSPEEDL@G���� �Ծ����)�9�����)��	)���SAM�WPx�0�1��MOVD�H$_S`Y%nk%$_��1�t�2�t�� ��c�v��8�H�PxIN����������(�+(+GA�MM<Vu!�$G#ETE�U�ٓD5��r=
�PLIBRv���]I�$HIu�_L�HݰpB�&E�(A�.� �&LW�-�&�,�)�	6�&1��f�`j��� �$PDCK����ٓ_���r �E���b7��a4���a9�� $I
��R�`D�c�b~���`LE�qkq���81�ƶ0���`Vp��P/aUR_SCR���A�r��S_SA�VE_D��8Ex�NO5�C��y�6�8@{$ E�.{I��G	{I�@�J �KP�q��H� ��� x"Mao���s� ���d��6W2U�Cqty� M� �k� F��aE��3�W<�@�[�jQWg@5r�U�R �R��Sc2jQM"��[�CL�W��M)ATr� � $PY��Ν�$W`�fNG �O�`�b�b� b#�HЈ��a� ���cJ��X�O���Z�e8��ހRt� p䠰p�3+zO�O�O�O�Ot�a5�_�r� |� E�8@��>vs�>v��8@�_�kwVvy�Eހu% Q��uB�\�P�"tP���PM&�Q}U5 � 8*��QCOU�1��QT�H#pHOL<�QH�YS��ESe�qU�E�p.BZ�O�� � q�P���%��UN\ְ�Q ��OE��p� P2�3��AÔ�ROG�����Q2(�O}�2�������INFO�q� �#�e����R��OI� (�0SLE�Q�с�рi���O�{�D��L��`� O�K0r��!E� N9U!��AUTTA�COPYqu�?��ъ`@ML�NI�M�X�C�ᐛ� Y�RGAD�J�q�i�X�Q���$ഖ�`��W��P����0�������EX�8�YC0b�O�bp�q���$�_NA9!�������`~��� � Q���POR�A�B��SRV0�)a�Y�DI��T_��{����Р���������5��6J��7��8y��S8BzL��m�MC_F�p
��PL9A8An�ȰR��9��Ѽ��$i�B����d� ,�0F1L-`L�C@YN�[��M��C?��PWR�c��L��!�DELiA��8Y5�AD�a���QSKIPN� �Q�4�OR`�NT�� ��P_ 4��ַ@lbYp� ���������Ƞ���ՠ��������9��1�J2R� L��� 4*�EXs TQ %����(Q����p������p���RDCf�S �`��X9�R�p������r��A$RGoEAR_� IOT�2FLG��vi��M%sPC��B�UM_��~��J2TH2N'��� 1�����G:8 T00 ����ЉMlѺ`I�8��R�EFr1�q� l<�h��ENAB{�(cTPE�0�1��� i�m���^QB#��:��"���� ��2�ҙ�����������&�3�Қ7�I�[�m���
&�4�қ��������(���&�5�Ҝ1�C��U�g�y���&�6�ҝ�����������&�7�Ҟ+=Oas�
&�8�ҟ����x�&�SMSK�q��|��a��E?A��P��MOTEF����a@��(Q�IOQ5�Ic(P���POW�0L�� ��pZ�����$�L���U�"$DSB_S�IGN�1)Q%���Cxl�(P�S232���b�iDEVIC�EUS�,R'RPA�RIT��D!OPB�IT`QY�OWCONTR;�(Q��O�'RCU� MDSUX/TASKT3N�p[0ހ$TATU`P���S�0L����p_�,PC9�$FRE?EFROMSp���%�GET�0�UP�D(�A�2��RSP|� J��� !)$USA^���6<���ERIO�P@&bpRY�5:"_>@ �qP}1�!�6WRKI�[D���6��aFR�IENDmQ�P$�UFw���0TOO�LFMY�t$L�ENGTH_VT�l�FIR�`-C�RSyEN ;IUFINR:]��RGI�1ӐOAITI��4GXӱlCI�FG2�7G1�0�Ѐ3�B�GPR� A��O_~ +0!�1R�EЀ�E3�e�TCp���Q�AV �G8��"J���u1~! ���J�8�%��%m� ��5�0G4�X �_0)�L|�T�3H@6��8���%r4E3GU�IW�P�W�R�TD�� ��T��а��Q�Tm�{$V 2���H�1���91�8�02�;2/k3�;3�:iva �9=i�aa�^S�jRS$V��SBV�EV'�(V�BK�����&c �p��F�"{�@�2q�kPS�E��$.r8RC��o$AŠFwCPR��Gv]U�cS'�p� 7�?8I�� 0�@DqV`��p�d`���PE0�@��=�
B5S!/� ��aRg�����R�6�N AX�!$�A�0L(A���r/THIC�1Y���h�t1TFEI��q�u�IF_CH�3�qI0�G�a�pG1bxf�з�m���S@��_J�F��PR�ֱ�S���Ԁ�d �$�SР�Z�GROU��̃TOT�t̃D;SP�JOG���#&��_P��"O������j��&KEP(�I�R����@M�R@�A	P�Qn�E^�`�!�[��SYS6��"[�PGu�BRK�B �.��pIq�p��M���΂��`AD�!̃9�BS�OC׆�NӕDU�MMY14�p@S}V�PDE_OP�#�SFSPD_OVR=���C����OR�CNm0�F�.����OV��SFR��pU���Fn��!#�p�C��A�"LCH�����РOV�s0��Wb�@M��ĥ:�RO�#�ߑ�_�p�� @�@�u@VER�ps0O�FSu@CV? �2WD6���2�ߑj2Y����TR�!���E_�FDOY�MB_CiM�D�B�BL�b>�f��attV"Q�240�/p��N�Gg�z�AM�x�Z�0���¿_M�~��"7����8$C�A�7�D����HcBK81��IO�5q���QPPAʀ=�"�M�5�͵���DVC_DBxC~� � 3"�Т�!��1�����3����pН�*���U�3��CAB ��2VӆPѣIP��c��O��UX�SUB'CPU�r	�S�P  P���90^SQ׹c��."~��$HW_C�А���S��cA�A�pl_$UNIT��l��ATTRI"���	��CYCL��NEC�A��J�FLTR_2_FI_�G(��9&��1LP�?�>�_S�CT�CF_��F_��6��FS8!����CHA�1�wᇲ�"v�RSD�4"�����q�_T��PROX��>�� EMy_ܠr��8d��a d���a��DIb0!�RAOILAC��9RM��CLOÐ C��Q*q���3q���PR��S�Q�pU�Cr�s 	��FUNC��@rRIN'PѸ0��u��!3RA��B ����8F�Ğ�WAR~���#BLQ����A��������DA����	����LD)0��Q1�q2��*q1TI2rQ�ǁ�p$xPRIA�1�"AFB�P�!�|ߠ�<`�R���MsOI��A�DF_&@؅�51��LM��FAށ@HRDY�4ORG6 H���A�0 �MULSE&@"�Q��a �G�	���m��$d$�1$1 ���0��߮� xm�EG0�̃�`ARހ���09�2o��z�A�XE�ROB�Wd�A��_�œSY������S�WRI�@s1��STR��� ��(�E�� !	%1��AB( �/&�a�ӰOT0v^�	$ߠARY�s�f"���S@	�FI���*�$LINK(���!�a_%#��%{q�"XYZp82�*�q�#OFF��R�"�"�(j Bဂj�4С��n�3FI��%7�q���j����_J���%��#�QO�P_>$H+5�3�PT�B\1�2C��i�D�U�&62�TURN��2r�5t!}��p��|7FL�`���m�0��%+*7�	� 1��. K�M�&8�2�Q�2rQ�#�ORQ ��G��-(�+p��z��� 3q�E"��T�GOV�@-A��M*�y�4 �E:�E@�FW�J� �G���D��o�*� � �A7�P��y��E�A�G`ZU:ZU�CG�ER�
��	6�E���B�TAFQ��)4����r'�AXУa2.q �c�W�c�W�c�W�p�Z �0�Z�0�Z%@�ZK@�Z ��Z
!�V� �Y� 
i � i� *i� :i� Ji � Zi� ji� zi�a�ioDEBU{�$v� u��;q��"F7O�n�CAB��6��CV�z� 
fr����u kњw�!�w�!�w�1�w �1�w%A�wKA�w��p\0��"3LAB"2�|EwЄ�҂�3 � EERVEN�� � $q�_�NAǁ!_�PO�����` f�M�_M�RA��� d r T���ERR��L��~ TYi��RI�qV"0�S��TOQ�T�)PL��T�Ѕ�-�����J � �p�PTl X���_VA1�b�Q���#�2�!2+�����/@��p��5�$W��V�����O�[�$�@�� ��S���Q�	EHE�LL_CFGN�� 5%�B_BAS��SRvp0�K� �S��JϐU1a�%Α2�3�U4�5�6�7�8�RO���� f� NL:�3ABn��АACKwv��)��o�u0iႩ_P�U2�COq��OU��P��ӕ������TP�_KAR��0��REm�� P8��z QUE٩����@���CSTOPI_ALzs��� �p��TĠ�� SEM[�dw�k�Mw�y�TY��3SO`��DI����p��=�װ_TMKӟMANRQζ� E���$KEYSWITCH��Ѱ���HE��BEAT4��R�EpLE����
&�U��Fd�����S_O_HOM� O��7REF�@PRi��R(� ��C@�O0�p �ECO���� _I�OCM�4M�k�pL���'�O� D�!$ۧH�U��;�M7�<�@�3FORCߣ�� ��OMq �� @Etxk�U�#Po1B�O�o3�B�4x_�SNP�X_AS��� 0�ݐADD��(�$�SIZߡ$VA�R�TIPr�q�G�A(ҷ��
�˨�r�t�n�SV�XC<����FRIF�R��aS%�7�x���NFѲ�EАO� x�PS�IڂTEC*�%CSKGL=�T�"�0&��V�D��>�STMTd
�o�P\�BW�@�?�SHOWw��P��SV� K�� ���A00�0�Q�� K���O���_���i���U5��6��7��8��9��A����6������20��F��
 �� ��U ����� ����0��� �J@��:�1G�1�T�1a�1n�1{�1���2��2��2��2���2��2�2�2� �2-�2:�2G�2�T�2a�2n�2{�2���3��3��3��3���3��3�3�3� �3-�3:�3G�3�T�3a�3n�3{�3���454��4��4���4��4�4�4� �4-�4:�4G�4�T�4a�4n�4{�4���555��5��5���5��5�5�5� �5-�5:�5G�5�T�5a�5n�5{�5���656��6��6���6��6�6�6� �6-�6:�6G�6�T�6a�6n�6{�6���757��7��7���7��7�7�7� �7-�7:�7G�7�T�7a�7n�7{�7ڈ���VP$�UP}D��  �Px���x�YSLO��� � ��հ�����QTAS�sTƠ���ALU}U����C�U��WFdQID_YLѳ�UHI�ZI�?$FILE_Σ�Tf�$u�_VSA��� h��+`E_B�LCK(�8bg�AhD_CPUQi��Qi����Sod_R1�ɢR ;��
PW,�d�[ �aLA�S��8�c�a�dRUN5��a �d�a�d��5��a�d�a��d �T�pACC����X -$&qLEN~�3t��&p䫠��Iѱ
�LOWo_AXI(�F1&q
�T2mwM��ɢ���I����Q�yTOR.�&p�{DW��s�LACE���&p�����_MAuйv�u�w�qTCV�|��wTڱ�;�1�<ѷt?�H_��s?�J����M��"��J����u���u2q2��������s6�pJKцVK~��4���3ՃJ0����JJ�JJ��AAAL�����4�5Xr;�N1B�N���	��tL�p_k���x@P"p��� `5`�GROU�PY�ӲB>$�NFLIC�ө�REQUIREv�EBUV�"q���кp2���#pɖ!qxг��� \��APP�RՐC���p
!�E�N�CLOz�,�SC_M ���A��u
!q޸�� 䣠MCp�r;�Xr|�_MG���C��,`��N��p��wBRK��NOL��t����Rϰ_LI��Hէ����JޠѤP� �p��p���p;��pD�"�p6�K��8�ц�>���� ҒMr�:ql�Gqz�PATHv�������Rx��������pCNR�CA���է���IN%rU�C�pwQ�Cd�UMB�Yop�����QE:p��Gp�����PAYwLOAͧJ2LHPOR_ANqQ�L�`�[�W�K�g���R_F�2LSHRё�L�O\�䱕����ACRL_�����޷�C�XrH�P"�$H����FLEX�� qJ%u� : 2Dv�p4�K�GYq�pPbt|F1Kљխ׀��������E ����/�A�S�e� w�����y���ф���� ������J�ÊT���X����υ ��څ�� [����
�� �)��@;�D�V�h�z���J��� � ��������QIPAT��ё��EML4� �ؘJ����ߐJE��CTR,ޱ��TN��F�ɗHAND_VBp�qѹP`�� $&��F2��K��ШRSW�b  qj��� '$$M��}�R��E@��Uw�H��sA�P H����Q���A���P
��A��Aɫ���j`���D��DɫP��G�`1)ST��9!��9!N̨DY�`���| �Y�鰋�KыǦ�J� ч�s�U�ХP�� &�/�8�A�J�S�=��� ; �t�.R66<N�/QASYM����	Ґ����Խ��ٿ_SH�����筈4@��+�=�O�JV���h�'CI����_V�I�dHN�u@V_�UNI�ÉD���J ҅�B�%�B�̦D�ųD �F�̓��������*UBc��ӆ��H�`f��XQEN� �v�DIɠS�OwT8*YP��� ��I�1A��äQ�`Bc��S`�  p�a.a� �� ME�����R'RDaTkPPT@�0) ���Qz�~����0�Xa	iT@�� $DUMMY}1��$PS_�гRF��)$Pf6�aLA��YP�jb��S$GLB_T >mU�e�PpQ p����Q� X	�ɗ`�SuT��ߐSBR���M21_V��8$_SV_ER��OÐL�c�cCL�`�bA5��O�RTPT O�P �� D �`OB���LO˰&uq9cp�`r�0�SYSq�ADR�TP�PTC}Hb � ,&����W_NA����tz�%�TSR~���l = ��M�u`�ys�u~ �s��s������� ����0�)�T�"� 5�~���B����s�?�?��?D��XSCRE�)�p�ȐST�[�s}�P!��tԈQr _� Aq� T	��`ob��a`�l�P�Ҥ��g�c�O� �IS�c��U w�UE�T� �ñ�jp^`Sq�RSM�_iqmUUNEXCcEPlV֑XPS_�a ����޳����޳R��COU�ҒS� [1�d�UE�tҘR|�b9�PROGM� {FL�$CU�`�PO?Q��*UI_��PH�� � 8\џ�_HEP������PRY ?���`Ab_�?dGb��OU}S�� � @�`~v$BUTT��RV`��COLUMx��U3�SERVx���PANE� q�:�P@GEU�<��F���q)$HELyPB�l2ETER��)_��m�Am���l� ��l�0l�0l�0Q�SINf��S@N0��� ǧ1����ޠ ��)�LNkr֓ ��`T�_B���s$H�b TEX��*��ja>�RELVB��DIP>�P�"�M�M3�?,i�0ðN��jae���USRVwIEWq� <�`��PU�PNFI<� ��FOCUP��7PRIa0m@`(Q���TRIPzqm��UNP�T� xf0��mUWARNlU���SRTOL�u����3�O�3OR�N3�RAU�6�T�K�vw�VI͑�U�� $V�PA�TH��V�CACH��LOG�נ�LI�M�B���xv��HwOST�r!�Rz��R<�OBOT�sV��IM�� gdS)�} 2����a���a��V�CPU_AVAIYLeb��EX��!W1N��=�>f1?e1?e�1 n�S��'�$BACKLAS���u�n���p�  �fPC�3�@$T�OOL�t$n�_J;MPd� ݽ��U�$SS�C6�QV�SHIF ��S�AP`V��tĐG�R+�^P�OSUR�W�P�RADI��P�_ cb���|a�Qzr|��LU�A$OUT?PUT_BMc�J�IM���2��=@zr��wTIL��SCOL���C����ҭ�Һ� ���������o�od!5�?��Ȧ2Ƣ��0�T���vyDJU�2��� �WAIT�U����n���%��N�E>u�YBO� �� $UP�vtfaSB�	TPE/�NEC��� �ؐ�`0�R6�(�Q���� ش�SBL�TM [��q��9p���.pv�OP��MASf�W_DO�rdATZp�D�J����Zp�D�ELAYng�JO ذ��q�3����v0`��vx��,d9pY_�р�	�7"\��цrP?� �QZABC�u� ��c"�ӛ�=
X`�$$C�������!X`�P<� � VIRT���/΢ ABSf�u�1 ��%� ?< �!�/ �/??0?B?T?f?x? �?�?�?�?�?�?�?O O,O>OPObOtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo Zolo~o�o�o�o�o�o��o�o{� ��AXL�MT�s��#  �tIN&8qtGPREO��+vup�XuLARMRECOV �)Xrzu�jF �%�!d�� ����7�I�[�m��~�,� �/��uN�G5� �+	 �A   ڏ�� PoPLIC5�?�%�upՁHa�ndlingTo�ol -� 
V�7.70P/36�뀬�
]�_SW�2�D�F0j�W� �43Y�J�9�K�7gDA7?����
&��X�e	-�Non%e��J����� �T7�	���E_�Viu�6s��UTOz"�,tTy.�?HGAPON� %���!.�U��D 1�y� t�x�����xy.�K�Q 1�{S  Hp�������	���uq��"=�" �!���Hեw��HTTHKY��"ٯ� ���u�����󿽿Ͽ �����)�;�M�_� qσϕ��Ϲ������� ��%�7�I�[�m�� ���ߵ���������� !�3�E�W�i�{���� ������������/� A�S�e�w��������� ������+=O as������ �'9K]o �������� /#/5/G/Y/k/}/�/ �/�/�/�/�/�/?? 1?C?U?g?y?�?�?�? �?�?�?�?	OO-O?O QOcOuO�O�O�O�O�O�O���TOĀ���DO_CLEAN�D���{SNM  ɋ���_�_�_�_o���_DSPDRY�R�_��HI!��]@ �_}o�o�o�o�o�o�o��o1CU��MAX �bTQNQS�sq�XbTB�o�B���PL�UGGb�cWo��P�RC4`B�P]k�lo^�rO�r=o��SEGF;�K�+�6� �_�_}�������ŏ�0�LAPZom�/�� +�=�O�a�s�������ໟ͟ߟ�6�TOT�AL�v�y6�USE+NUZ�g� HXL��NR��RG_STR�ING 13�
_�M,�S��
��_ITEM1��  n󝬯�� Я�����*�<�N� `�r���������̿޿���I/O �SIGNAL���Tryout �Mode��In�pB�Simula�ted��Out�T�OVERR~W` = 100���In cycl�Hŕ�Prog OAbor^Õ�>ĿStatus��	�Heartbea�t��MH Fa�ul����Aler �����'�9�K�]�po߁ߓߥ� ^S ��^Q��������,� >�P�b�t����� ��������(�:���WOR9���r���L� ������������ *<N`r���p����PO�� �����9K]o �������� /#/5/G/Y/k/}/�/DEV� -�/ �/�/??)?;?M?_? q?�?�?�?�?�?�?�?�OO%O7OPALT��^A��8O�O�O�O �O�O�O�O__(_:_ L_^_p_�_�_�_�_�_LOGRIxp��avO �_*o<oNo`oro�o�o �o�o�o�o�o&@8J\n�_*�R�� �qo������ (�:�L�^�p����������ʏ܏� ���PREGbNK��$�r� ��������̟ޟ�� �&�8�J�\�n������������$ARG�_r�D ?	�������  	$�W	[�]����.��SBN_CONFIG ���L�K�F�CII�_SAVE  ��k�b��TCE�LLSETUP ���%  OM�E_IO��%MOV_H��¿ȿ�REP�|��UT�OBACK���V�FRA:\8� �8����'`��8�c�,�I�NIa@8�^�~,�MESSAGz��������ODE_!D��}�C���O� ���,�PAUS!�~�� ((O�� J�\�F�|�jߠߎ��� ����������B�0��f�t�%�*TSK � 5ݒϕ�/�UP3DT����d�����XSCRDCFG� 1��� 	�������&�8�J� \�n���\�n������ ����"��F��j |����/e�>2�GROUN��߾�UP_NAܰ���	2��_ED���1
��
 �%�-BCKEDT�-��}��pDg�Ӱ-2�p8�/�Y/�8���g2���E/��/��/8~/��ED3n/&/��/J/\.�/"?�/�/ED4?�/?�/\.[?8�?5?G?ED5�?n?�#O�?\.�?jO�?�?ED6ZOO�O6O\.�O8_}O�OED7�O�O�k_�O\.G_�_!_3_ECD8�_�o�]-p�_Vo�_�_ED9Fo�_�o"o]-�o�oio{oCRoY_Vh�]�1�{� LNO�_DELGE?_UNUSE	�LAL_OUT �V��WD_ABOR���~�5�ITR_RTN��=�H�NONS)Ю������CAM_PARAM 1�����
 8
SO�NY XC-56� 2345678�90Y �f�@����?�W�( �А��8�h�х�:ڎ��HR5ǃ�ɜ	��R570�B�Affފ������ ڟ�ǟ�"���F�X��3�|���i���į!�CE_RIA_I�������F���;�Я ���GPw 1��A�s�����V�C�Ҹ�����CO�C ���(��ǀC8��@2��H��CCX�����Ch��p��x����� C������ ���+�=�G��ށ���HE/pONFIG�=�f�G_PRI 1�B�$r�π��������(�~�C�HKPAUS�� 91���� ,wuj� |ߎߠ߲��������� ��0�B�T�f�x��h���D�O����T��_MORGRoP 2?� �\�� 	 �,���P�>�t�b���5���H��e�.�?a�a�����K���d�P�|V��a�-`�/A�

s��@�����b&�i��.ܦPDB������)
mc:cpm�idbg��:_�  �+�����p�U   ��_ ߀
�3�� ��d����r}C�e�*/��/��{g�+/$�g��}f/s/�i�u/�
DEF ��(K�)�b b?uf.txt�/\�/��_MC����E�d,53������ʇ�Cz  B��p�B�Z�B��X�B��~B����B��C3��
q�Dv���D:�"Df���DRt�DG}S�D�a��=F�p�gF=C�Fi��WF�EF�2�?FjI�	ބt	6����4���(D~���/��ʄ3@à1/�  TB�D.Da�  EI�5� �F*� F�G$�ˀF[� GR��kNGl��G���G��&H���G֓�H���߃]��  >�?33 �ށ��  n^��@߂5�Y�Ed��A��=�L��<#�
 ���_�*2RS/MOFS��.^��9T1��DE ���l 
 Q�;�P  0_*_>/TEST�"__��ER���#o^6C@A�KY��Qo2I��B�0�� �C�q�eT�pFPROG %�S�o�g�I�qRu����dKEY_TBL  6���y� �	
��� !"#$�%&'()*+,�-./01��:;�<=>?@ABC�� GHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾�����q���͓��������������������������������������������������?������Eъ`�LCK�l���`�`S�TAT�c_AU_TO_DO���O�INDT_EN�B;���R�QY�K�T92����STO�~���TRL�`LET�E�ފ_SCR�EEN jkcsc 	��UπMMENU �1i  <�l�ol�K�u��� FS����柽�ϟ�� �R�)�;�a���q��� Я�����ݯ��N� %�7���[�m������� ɿ�ٿ�8��!�n� E�W�}϶ύϟ����� ��"����1�j�A�S� ��w߉��߭߿���� ���T�+�=��a�s� �����������>� �'�M���]�o����� ��������:#�p)+�_MANU�ALӏ��DBCO�u�RIG�$�DB�NUMLIM��,1e
�PXWO_RK 1k�_�-<_N`r�T;B_�  m���Y0�_AWAYJ��1G�@b=�P�_AL� =����YҀ��`�_�  �1!�[ , 

:&d2/o/�&�%Mt�IZP�@P�#�ONTIM��&d��&�
�e#MOTNEND�o�$RECORD �1'kU2)?�!�O�?1-?&k�k?}? �?�?88�?�???�?c? O*O<O�?�?rO�?�O O�O�O�O�O�O_�O 8_�O\_n_�_�__�_ %_�_I_�_o"o4o�_ Xo�_|o�_�o�o�o�o Eo�oio�oBTf x�o��/�� ���>�)�7�t��  pu�����-��͏ۏ �����N�`�Ϗ��o� ���)�;������ 8���\�˟ݟ����;� Q�گI���m��4�F��X��TOLER7ENC�B�	"��L�Ͱ CS_C�FG ( +x'd�MC:\��L�%04d.CSVdY� cֿx#A ��+CH�z _/x.��G��},��RC_�OUT )��- z/��SGN �*��"��#��08-JUN-�25 13:41���27-M{AY��4:38��]� Z�t������x.����pa��m��PJP���k�VERSIO�N ��V�2.0.11~+E�FLOGIC 1�+� 	d���ٓ��p�PROG_ENB�2��WULS�' �p�_WRSTJN� ���"�EMO_O�PT_SL ?	��]�
 	Rg575x#?�74D�56E�7E�50i�dԂo�2E�d��j�"�TO  .����k�[V_� EX�d�%� �PATH A��A\��M�_��~+ICT�F��, '�`��eg��}�STBF_TTS�(�	��E��`���� MAU���ߧ"MSW��-D )��},t���.�!��]l�R�v������4SBL__FAULy�/�|�#GPMSK��^�"TDIA��0����`���!1�234567890xS�l�P��� ��//%/7/I/[/ m//�/�/�/�/�/LZ0PV �� �/�2?X?j?|? �?�?�?�?�?�?�?O�O0OBOTOfO8<x�U3MP$�I� �A�TR>�O�@PM�E���OY_TEM=P��È�3��4󜐰�DUNI	�w�Y�N_BRK 1���x�EMGDI_�STA	��_�LPN�C2_SCR 27[��_�_�_�_ �&�_�_o o2or�nSUQ13y_+?|o�o�oвolRTd47[�Q��o�o���_>P bt������ ���(�:�L�^�p� ������ ?Ǐُ�0� ,p��+�=�O�a�s� ��������͟ߟ�� �'�9�K�]�o����� ����ɯ�����#� 5�G�Y�k�}������� ſ׿�����1�C� U�g�yϋϝ�ׯ���� ����	��-�?�Q�c� u߇ߙ߽߫������� ��)�;�M�_�q�� �ϧ���������� %�7�I�[�m������ ����������!3 EW��{���� ���/AS ew������ �//+/=/wa/s/ �/�/�/�/�/�/�/? ?'?9?K?]?o?�?�? �?�?�?�?�?�?OK/ 5OGOYOkO}O�O�O�O �O�O�O�O__1_C_�U_g_y_�_�_�_�gE�TMODE 15v'Efa t�|�_GgRROR�_PROG %��Z%���HogTA�BLE  �[�1O�o�o�o�ZRRSEV_NUM �R  ��Q��`a_AUTO_?ENB  u�S�Zd_NO�a 6��[�Q�b  *U�6p�6p�6p�6p��`+5pOastH�IS�cXa�P{_A�LM 17�[ e���6|6`+t����&�8�J�x_\�bp  �[4q��R���PTCP_V_ER !�Z!6o�Z�$EXTLOGo_REQ�v�y��SIZ�܄TOoL  XaDz�r��A ܄_BW�Do�%��fQ���_D�I?� 8'E�t�TXa b[�STE�Pg�y��P��OP_�DO�v$v`FE�ATURE 9�'EQ��QH�andlingT�ool � DE�R Engl�ish Dict�ionary�7� (RAA �Vis"� Mas�ter���
T�E0�nalog �I/O��p1�
0�uto So�ftware U�pdateb� "�/�k�matic �Backup
�d�
!��gr�ound Edi�tB�  25L�CamerazT�FX� "Lo���ellT��L, �P��omm9�sh�ۡ�h600��c9ou���uct��p��pane� DI�F���tyle �selectѡ-� /�Con��9�o�nitor��H�d�tr�Reli�abT�ϣ(R-�Diagnos���Q�	�H�Dual� Check S�afety UI�Fc�Enhanc�ed Rob S�erv��q ��v	ԸUser sFr���T_i��xt. DIO Vf�fi�� )�\�wendܰErru�=L��  prנ*��rO�� @���EN�FCTN M�enuİv����.�fd`�TP In�?�faco�  
�E�G��p;�k E�xcذg�C��High-Speܰ�Ski��  Pa�r+�H���mmuwnic��ons��7\ap��urf�?�~X�t\h8U�^��connZ�2Т{ !�Incr���str)�8��M-�6�KAREL �Cmd. L��u�a��}��B�Runw-Ti�Env��(<�@�I�<�+��s���S/W�"H��License̾��� ad���ogBook(Sy>��m)	���"M�ACROs,��/_Offse\�f��b��H�!�Y�M1��MechStop� ProtZ�3� �5
�Mi4�S�hif\��B6S�MixܰQ�����H�Mode SwoitchY�Mok�*��.�� ��Mt�Q��g�� �5��ulti-T������)��Posj�Regi�>���  ! �P>A�t Fun1���6iB/��R�Nu!m�Y�3�G�P/��>� Adju��	��/2HS�)� o<(�8�tatu���wAD ��RDMޱ�ot�scove&� #e�v�㱗���uest 867�.��o�\���SNPX b��Y���)��Libr%�
�rt I���� "�����.S�o� ��s i?n VCCM����� j���������/I�� 710~�TMILIBXp����g�Acc��C/2�TPTyX�� �Teln���Y@����K�PC�Unexcep�tܰmotn�� �������\m725����w�5����  h640SP CSXC�i � xj*�� RIN��sWe���50,��vrl�زmenX" ��fiP-�a��x�P��Grid{��play F O`/��? ��ELR;��|�20��ORD�K�sciiw�lo�ad�41d�st��Patd��CyqcT�h���oriɰz:�7c Data� qu6�2�0�*��������FRLa�mc�K�HMI D�e��(����k�PC��φ�Passwo�rd�644��S�p�����D#YEL?LOW BO�	?1��Arc%�vishu����#ti�Op��^�! 2��aO�p�o�� t��ֶT1�o�����HT��xyy�	�   $�t۠ig��10Ơ� 41\+�JPN� ARCPSU �PR+�8b!OL�0Sup�2fil�� �!��E@-�;�croc�82��v���$� 12jSS0e.4�tex-� I�7��So��tf�ssaEg�� e��У�P���,��� "Tc Vi#rt��v�!����gdpn�
�J3��SHADf0MOV�E T�MOS �O TԠge�t_var fails l�>PU~1�E���� Hold_ Bus %�h���VIS UPDA�TE IRTORCHMA A�{�vY�WELDTV S �]�DtS: R74-1��ouiPb}�y���BACKGRO�UND EDIT� "RC$REPTC�D CAN CR�ASH FRVR� 62z1�SCra���s 2-D��r� ) "��$FN�O NOT RE���RED �` m� ��JO� QU�ICKaPOP FLEN m41S��Loc��gRTIM�Q%�#�FPLN:� FG��pl m�r�`�MD DEVI�CE ASSER�T WIT PC�V;PB�AN#aAC�CESS M .�pc��Jo��Quqi±�Kbldmg�USB$ ��t &� remov�� �Pg�SMB NUqL� ;a|�FIX��}C��ACHIN,Q�OL�`MO OP�T ՠa��PPO�ST0�WDU C��wQAdd�`ad����0io�2��$�P�`W\0.$0`O��IN&�P:fi�x CPMO-0�46 issue�C�J/aO-�0�r1�30Т- ��vRS�ET VARIA�BLES-P{��R3�D m��view� d��M��&�ea����b��of F�D�5P:N@x O�S-1y0`�h s�c���t��s t�l�o��7 WA�PZ�3 CNT0 T��/"�ImR�)�ca� �Pu��POT:oWhenapewB�OSTY E�{1t���ptKQdo GE�T_�p �p��VM�GR LOl�REAd0C~QW�~1�(�pl�s�gD�ECTp�LpING IM�PR�DR(p+PB�P�ROGRAM�ER�IPE:STAR{TU� AIN-;��ӠM/ASCII<zPÂOF Lq�DPTTB: N�p;ML$me P����`:x�mo&�alqlW`!�ӤTorc�!A�U�HC�iLpԸ�th�`n�@ ch��/GEA�!�tou<͐�RCal��k�oSign`� ND��ԗThresh1�23��`��09p :? MSG_P�+0Ger  �Q�Aܠ�zeron��0 gH85��RImA��n�2D��rc�0I���OMEa`�pON�aP5�  נSRE#G:FF-Д� ]�'����KANJI��nʖ�J��c�0asn yd�!OA immc ��INISITA?LIZATI�����~1wem����dr>+� LB A�UWq�minim�reAc[�c!�R���m$�ro -1>ѮS�ܰir��@ұJ�1pd�ETw�� 5`?�I�o�w u��< se W1lc��YbPM����p�Q���R`vR&�lyu\�3�Re 0�d4q�q1#���m <a��arn��ঁB�ox fo��*PR'WRI�PW�S��v�k09 F�pupᐿde-rel2 d��p� j��`━be�twe��IND �Q���igE sn�ap|�us��sp�o TME��TP�D#�DO�p#aHANDL 1\k�`(vR��ȀD�ny�S��v�Yoperab�il� �T*�: H$ � l\p��Vq�b��R�< p�a*�c&2OƝ`FA,�.�-QV7�. f.v��GT�pi�s��� ɠ�tmLine-?Remark ��/ RM-�` W�#SPATH SA+P�LOOS UIF�c�+5f fig�pG#LA����Vrp����z��U�0ther�>V� Trac���tW�\b�s7��d�ht�� n�@  ��R�3:���dK�y���it k8�d�Pa�yR![2]�ü1�: g��s��doew�XQ��0IS�q��qEMCHK E�XCE C���M�F +�Xah�� 35\k��)���QBt���'b���[�c���e �`k�S�� BUGr��cD$`PETp����f�c4��0XPAN;SI��DIG��@�OoPmetTCCR�G EN��CEM�ENT�A M̀K� {�`H GUN�CHG �`� EX�T�P�2�bQS�9�3 wP8�x�ORY�LEAKq  H�5gyq�PLC W�RDN R �O �/u�QSPE=p��G*�V ��$�tn7w20\3pGRI���A�rT�PMC gETH��pSU7p��`  j5/n�PENS�PN,��*P� ont�`BRO�W�`!sRMV A�DDz CN qD�C���PT3 AL�A2@ ���pSVGN EARLY�R��ŰH57�Ga�JLAYҀE (�@M�PPD�p*@HΐS I`P�OU#CH8���V�F�q��comH�x ��ER�ROR� DE n�J��RO�CUR)S8pI��N4q��-158n7�R'SR xP#aUp��(�Rqy�T�Fz�;`�pk��t�� gՂ��B�SY RU;NN�  a�`��BRKCT�!RO<�p3@ \apSТ�cAXxP���h8+ <q��ISSUr} �sPX�PTSI�K�1M10_�IPSAFETY Ck�ECK[��Á�������<#X�� �TW�D2�@�@�INV���D ZOp�5Xx��t�DUALy�� "M6�0�"rF�#�E��dPdNDEX F�t*UF�"Pʀ�0sF�RVO117 A��PT6�KtqFAL�PTP2477D6r_�P�!;HIG� �CC�t;SNPX� MM��tq�d~ҁVq�q#�
"��DETEC�Tq*@RRU�qA�P�5p�9� y�)<9���7T���Pds� k��	���!Q���� �t\4A�;A0�2 "Ke@" 8@HI�q�XF8@4@H�PRDC"�
�aMB8@�IXF�b���zOX@8@���a�G}E�B�Ccscr��J8@�Ndctrl�d.�A�NZE�A5�$�Q��!�`�Df8@�`�m�878�Q-;� ^��� rm`�
���PR̠78�@RI08@0q�Q (~\Mp@��0t��!{B8@\tQ�<OX�St0�3hB3�nO�Vtp�A�@LC�F�L��� �Rpl�cf���J8@�WTam�ai�E8@mubov 2_miTA�O�S8@U`T[xtT�AqPr674xS�Shape GeQn��8@j�I�[R�`ĝ@8@T����%q (u8@��II�^�Q~C`�a�[8@;Ynrsg0��4� � 4�CtMr)68@�r5hB5�zVnnretsp "r��Po�wng0bGC�RE�Ka�ޠ�D�AT�E�k�creGat.�q�M�a�o|ksqgtpad1P<��(�tputZj�{ �������܆28@��0��Q����sl�o��;� �hexH�TBp�8�ď�keyH��8@�pmZb�NR�u7A+�nrgc8@UQ��pp�bUZ�dp0aj9�21xSpl.Co�llأcq�\A��RN�q�UA� (J�8@ip�_�WA��_�Y��ae7hB7�ͦtp[�? "TCLS9oKb��clskyh[��s�pkckZd����$�TQ���dA�rx�7�10a- KARE�L Use Sp��FCTN9�a�70l�0s0a�� (���a���~C8@��MI��c8�hB8"   ��8@ v	��v	   lm7atea99�qM�����E�mcclm5�CLM;�� �j��fE�et���aLM	��h�yasp,���mc_mot�B�N��8@0H����Q��su'��Q��ȕ�䅮���joi�#�ߕ��A_log8�Z���trc�B����ve�ϓ�v��QWX���6�finder�xSCenter qF1�lSw520���ha6rX� (<�r,�Q�Ձfi�Q �NH 0�I�ۡ���A8@uL���tq�a "FND�RVϳ���etgu;id�UID�C8@����������TA@�nuf;��P���ƞC�B��_z�Ӡo��qG�������l���fnd�rTY��2䁴tcp<"�,qCP MF�}�38@517��6s38�E��gf6��(� �K��Q��-�X��A�tm6�P�İ� �Q���	�͘��Ctm�Ĵ�b8@ej��TAiex��aP�Apa�ذ�cprm�A���l�_vars ��
��dwc7 TS���/�6��ma7AF�G�roup| sk ExchangJ �8@�VMASK H�5�0H593 H�0aH5@� 6� 5�8�!9�!8\�!4�!2���"(�/��;OMI� `@a0hB0`�ՁU4U1#SK(�x2�Q�0I�h��)�m�q�bWzR�Dis�playImQ@v�J40�Q8aJ�!(�P��;� 0a��0���� 40;�qvl? "DQVL�D���qvBXa`�uGHq�O|sC��avrdq�O�xEsim�K40sJ#st]��uDdX@TRgOyB�Bv40)�wA~����E�Easy N�ormal Ut�il(in�K�1?1 J553m�0bD2v�Q(lV40xU)��������k986�#8Uϕ�|�rP "NOR��dw d.a}oKksu�O�W���OY��W`�j0�6�H� me'nuuyP6�M�`wR�X�R577V�90� �RJ989}�4�9b\�`(�fity�����e�<?��&Vsmh`��8��C0�Sv�q�8���w��pn "MHMN <��ޣx�Ay`�o�3�u �`f�І�x�t��t�RzQ��LV��vP�tm����|I�1{oPx �2�|���I�3I/B�od3stǏًmn���^�}ensu_�L<����h!!��Rt��huserp��0Ҹ�ʐcM�_l�xP�oe�<�рpoper���>�xdetbo/�l> �x���Ps$p�`����OPydspweb ͓��z'R��u�Rr�101&S՟{t�`2�Z4�30�����"�`4�
�4�5��KQp�m[T��dUCalG 40`�Q)p40}������9;��DA�� �v	LATAum�pd�\bbk96M8��68c�fbl�.41969y�9�|�D����bd� "BB�OXêM��sch�ed����m�setauM:�����ff� ��40��n�41�ϒ�40�q�col��|�1�x1c�ؘ���li��X� 0���j��&�8�4 <�{ro5�TP E�l#��ryK42r���;�(T+Q �Rec'�ʈ1Iw�84��x���Ak971���71�;���parecjo��QNS��[T���dXrail| nagek�M ,QjT2 *� (�ĜR%<x�80!bTh��p��4��4�y�Dgl�paxrmr "XRM�g�l��brf{���n��k�l��9turbsp���㧑- �l015	�g�625C�Mh� +���)89��	+��B6��o�ҹ��x��7�q40����pd? "TSPD�=��tsgl��l�:`dQ���8Bct���K�vrE�aܮ������  1�!���21�`( AAVM �2��0 �@fd T�UP him (�J545 ly)�`8 616 %�VCAM ��CLIO (��0:�5&  (=F\ MSC �Rt"�PBsSTYL��D!28 :2\ N�RE F2h SCH�6pDCSU� tpsh �ORSR �rD!0�4�SEIOC�& \fxh 542� LEX"� ES�ETn�8!H ��sh�8 7H �MA�SK�Ø"7>��OKCO*`x�!03"6(�!/400:66$ G6s39.6[8LCH!6oOPLGR703
5OMHCR��0C� h(! �06�A.f8!�54
��00DSWb 588�180 �h!�37 88 (D��"02C24���27 q9�25��2-6��05��9PR�ST bBFR�DMES�!zB�9�30 _ NBA�  6� HLB �3 (~!SM�@ �Con� SPVC� �8!20z��T�CP aram\TMIL A���@PACETPT�X �@p TELON 96��29�%�UECK��r U?FRM et�P!�OR ORP IPL^%CSXC�0j�1�CVVF l F�QHTTP st�A")�I#� CGHP8~ZIGUI�0��hPPGS To�ol� H8�@dj`Z��!@�h!63�%j�@32Q\�31 B��h!96�%R651��Rs�!53 TF�AD�R41�8"1� ��oo�"9��41775�"/@�P�VCTO�@�U�!sh!{80�%PRXY�R��!770 �b8 8�85 ol3P� L� аdi� �`ڳh �LCP{Q� TSS� �b�26:����@C�PE �HT@VRqC~�tQNL ��@002 %��b	0gdis� �`7 <°�a\0�T�`1 �`e=n�b4 652�`)FU02Q0Πo`p2�Ptu�r4 $r�5N��RU0p@ns�e�QJp1 APFiI[ Jp3�g34�g40 alxrE1�t44w46� ts U0  7v�0O��r5�e�p7 p 7"sw�a61:��rY4��r5 QpwGr�`�$�p8R�"sP`tjQ�b�36w77�wL8`�v83���r8�&�:��pOq8�8 "r�key8�9F��a90�91 p�#@���� �D095�g97*pur�A1@d��H�P|P�q1�0QplSqA1p#4��]a!s1@sl༂8�Ӽ�\1�d1�`��v�@{��14p�ae��5 hH2��`�6ޣ��7�f1p@��d�YpCqd�ـ
d�1�`uq��� Cu�1< Oq� ��7ReU	1$ �u1�Pϱ� ���@- WQ158� ase C��9� B��60 82�ń�p���4 (W�ai��`吢!��7�E��8�EU1P`rIo9�<�1��<�2��<�	0��T��l�5HJ�l��cC���9%�GMCR��P�2�`t�Q2@967�QR��8��9Z�2TP�B���P�2P7U5 @�o���
�5�`U���3 w���?A�E$�1��c�qAwl��A��1��512 f���1�u5Р���a5p$��56�+a��Q15h��Ұ�1 @���pp�b[�538 BxaB��|p�4�2�1e1/q5�p�4U5�P16 (߲�Pz��0��8�P�����p�e5`�e5(�/�P`bbf>�X��$Z�U�}5d�\� X¿7 	  ��8� k_kv��79� s�82 &�H�5��E6���p����h ���ñ���3J"�`n��4 3Ȥ59ѧ�6�0t���8��6�D0$�$�4 7���!���<�j670\tchk<�Ps��<�B<�90��7�<�$��<�\K�<�q�Ӻ� A�C<���q�<���<�mt��sg<�lc���FA<�H��<���0<Я���<�hk��<� ��B<е�o�<���<�x�K�<�dflr��<Ш��� ��o�`����D�;�<�gEvam����B<г�oќ����<а�KЀ�creexl����P��<�X��|���j6<�s��prs.`���\����<�7������fs�gn��P�b�t�at ��<�L��1B !��svsch/  �S�ervo S��usle>�SVS��44�1u�_<��� y(����ched���,��~��A\��  �� B���B�qA����Zcj�� � 5��1<���Ә�p�cs?s "ACS<�& (��6� �����c el���Q����?torchms�<�7- T�Ma`Ѵ���09 J5;598 J681s�7� 8��b��<�p�a����te,s������/�E�� �m��ARC.�� 1q�4�!=��C�tc�pA�@t��Ѧf� F����7#�2x�SE�r���UstmS�0960'���RC����0��� p��96G= '��"H5W����L���\f�� �@PATb���`!4U�#!Stmt�E `��� �pMA�!�p��z�2?�in_�<�X��r�X e/c�W����V����e�tdl�vߏ\ov�eto���܏��m?monitr�\��|#�0st��?.6�a��PP���!� Q�!y`�`ame� �Arol�c�43�0 �p��ћ01� 25� � �<� v�	�v	�A@�818\n; <s�I��B�2�pMPTP"���C�1mocol ��,��CT�v�'!� �A����8P53��y`T/ouchs�s�`��<��J5���Ѩ`mP����n[PQ�a ,�E�a��IP&
�Pth�A<�KF#R�m;ޱQetth�TH�SR'�q-�Rt��o? "PGIO�#!$�s�ISwka�"WK���!�MHqH5�4��5w5n/�Sm/��@ 7�*�da���8`!w/Ac��tsnf Tk�/�#gb�aP��u`��^m�`u��Zӭ�ܱQp�є�#����Ka<��M��t5 QtZ�a<��dFS5GhK����G�1or��dW��64��tPx���P ����x,��?�$���P<�Z4e7�g? "SVGN.ox��copy "CO�;�Wj$�O�A�9� "FSG�ѧ�%7��_j��f� wQSWF*|!"(�sgatuɀ����_
��tp_T�PDo��9�79��#dߎ?���h�GA�T���!#��  �Гf�` ��"/� �w�Z� �b?6?� � ���� ���E ���M� �chrT� �K6K� �sms� �o6�ѐ�?gtdmen?3 ��?��� ���mkpd�td2 ���, ���pdQ�X� ����� ���mvbkup. ��[�C�С��mkun�o��prp���mk�l �4��s �nixU��� �ldvrw���glg�4�� ��渣���aut7�.pб�旐 �ַ������su3� �Ǜ� ��Ƿ� ���\ �6�b2X� ��&�� ������A4�  ��B   946" ���fB� �t\pai�c\p4k947� ���F#���� �icgtas���pa`���cc:�<��o���N��gen�� � �F�lnp � ����sctf@��1��wbO��c��Ջ�`��߄�vri�ߢ�а�-T� �x��p�flow� 6OPAc��ow���R50qtS �#T� (A��4�#���p��V�cu3�QF� �̾SI�ac����46`����s&��pa��`!!���� ���55�b  �o)�p���0娿
��afcal3�P� @��f��}���`�f��m	߳�p�d�m�/���a/��$C`ѷ�� �! track\P�� 0�ine/Rail Tr�]TJ�s69W�T  (L�� 8(`љT.�`�%��HD��P0� (��8��48��_ɛ�⇒4������ �3�b3����alV@ �N�Tf���%��Iinp]0m���aen�� ����&?5�c@Itst3@��$�� ��`�,R9�%���0�氱%��pope/ners-OW dGDev��F�M�6W����|A�Pc"�l!esv� �,��R��V$�Q`���U<�V$ �k9j 
�6��# �����%�paop/!OPN�U�V ��2celL��8g_��/�6��tscG��$��V!��3� 5vrop�ߡ�7`�n(`�V" 2D�a V'O$:S9�>�� PumpE�� jQ�@�" ��!
��@бMSC#�@��)P��AC��`��� � v����� \mhplug�@g�"7P���uK")㠱io7�CpJ0��E�LIO q51g 7A93շ�E5 q9 t����4rb� ST��R��CPJ�989�P�LSE(�' �e C3Q(P �/Ov���o�P�� ? I1�R���55���f�I1`�tcmio��MIO�����U�tco1"CL01dV �cBK`io��uM?���Sl�I0�߈��Eg �o���f �tI4\onfdtI����e%�p27�Inte\�TB CoMoo1�E�R�(do55G4 (;r>Ex,�8�nR##ipc�/>�&�qp5���
oQé�1�p����7/o���r5a�pd�CDV_���rP�֮��qp2cnQd��s �p��a�o��r`҄�S��"�c�a�c���2kIԿ?A�pcrt���or0�qd#��"���3p+����D��Џ��vr2k �0���AG�.+��gcho�;�uC��8(� �uV630�fw e P�mී�@���`���TX�� ��d�chp "_��(	��3�����8����\p3�v����ш�9��3�1 �����laow�[ͧ���chk���㳦s��s?Ө0�i�1h���2��i�w����s?1*�-	�:�O��vr������p0�'���PFRAPwWat?1rneE� P�sp�& ac5� _A.�rbo#�,�a��g��������Qs<�ICSP+ 9�_����� ���F�A9PH51IQ9%3 7��HX6hQ]PdVR`S5��fPR6 liQWPR� (P!/am S�u�"�A|�I0�tpprg�0���`h�@2atk932�!��E�^��a/sc "8�C��S>i�atp�"�d�@1�I�
g�dsbl�fltJA�Qsab?le Fau�P{�C!��EV0ex/!D�SB (DC��t �$�p��X 7� �� 5��Q�t3*�~��6��td9� "!%�(5��sb9኏����\	�6#���@5�p$�D@550-Adj�ust Poin	tO"tVJ�Rs�z�� ���!�X_�Yj��/0\sg��4��}7�y�\ada�"A�DJ���j�Qet�sha<�SHAP8�sŭ'jpo�r4� t�!��$ ��C|��	Tk!bRPKA�R/Qiagnos�tì!O!vV66C J`ew0�(��L���/�&krlde� ��PP���hUH b���r3�Pp?q���DBG2C��� ��X�o�1U�� `��WT`�@ipJC�M�aipper �Opv`1Se}78? (MH GF�  ;":�&##�� a�x��,�$��388C���(��#��9.�9C��g$##PPk�Q��8�!�_ "$�"��=0%�P��A $���_�#%0AQ�C~2 �Mat.Hand�lE��!= &�pq M�PLGET�0�1( �3�Tt&P�Sٰ'�B� 1��B0����&p��H�� PP �'p��@�C7PP@	�TG�tD5�}m�q��Afhnd "F~_R  �����>PP	   xT?Qܣ��P(Pa��To������?�pmpa�O��JP ak925B��2`@O�JRpsQ�`B2�unLHP�Tgse�GSo1�O�W��QT��v !�R�Pt�p~���JRdmon0.�@��V�!ns�hYvr�QJ�g�Q�o�jXY�HS~7sl�f ��pen�PDnR(R&���ɐ823'��ٔ q���g� ���� 1��� S�� ? �c\sl tQ�!|QE�P��a�rtP�g��P�� �v��"S�EDG8�s0�qtdgY T����v P`ho�s`<`����qc�`g
�e` o�w8�a@o"�ile6�H�e�ȅnR�� �e<! j517�>����J%��e�`��BQ4��Q&�L�!F�J�=�o�5�z/l17���_�œ��`C�0C�  ���LANG j��A��������gad���,#�jp�.��4�Ē�ib���s�Ƒpa���&�~��j539.f��,Ru� Env�
������3H�z�J9�����h�Ф
Ҕ���2�2����� (KL�n-TimФ�⠤���p�3�TS����\k}l�UTIL"o����x�r "QMG�l��!������1 �"��S�T3�\kcmno��SФT2�椱ut�.�lre3adc�}�exY�ܤ�r��\��l��Фw�a3��2C�*� -� C�D�E!Ĥ� .��C�� R CV̴�Ҁ�\�p�Р���p�t�box��.�@�cyscsL�:�RBTE��veriOP�TNE���;ӕ�k�e`�ߦ�a�ߦ�hg����DPN��gp.�v��r�ptli�t��0�4��te�\cy����tmnu3`�r���5UPDT��������駣��it�e �� swtox�,���oolB� F"�Y���Q��(q��gr3��䪒��"�䂴�w������߳��s �������������ylS���bx "O�� ����l����P���A�l\t�� ��p������	�Col�9e!��R C��r���&r �m;`��Chang�Lq�T1 �rcm3�"��
� A6���"����sP7���"��222���2D45�7�� CCFM��H��accda��Q�c' ��KÕ 0���K!����mo!�� �,$Á��!"
� ���/�/����	Y�,$0��)�,$sk����
m rC%tS1,$+��<k1�%unc.,$o�8��1��sub����8��1��cce�5/�!&��-/?-W/i&v s�}/�%#�#�/�.C� �/� C%
�@? U �&�+��F:qt�
pD��� D	  �U�:7�Dxmov.�P��DPvc5Q�tfr@PeC_UYg�eobdtg_y[tAu���P���PTUt�P��Sx�_�^z�_�\v3ar�_�\xy�_�[pcl`c�P���P��Ue�Pgrips9uaoskuti���o>vfinfpo}��o��j�b�P���Qud\@�aX��Pc�\Rrp�QAnƅ�P�v�P)tm#q`Ɔ�P�v�a+rog�aࣆ\Q�?a+rpal?a{�{spa���P�u�Q�t�_TZp�0�osi�pkag3r�ovlclay(�:�t�p�T�d�pu?a�c�A� �����KtKa�P����9qTf|rdm��{Grin#r���s� �2���|s�Pd�v�tv��v�h�0��yGstn* џ�yt'�	1�p��D�p�uϑ#�Cul�@o�W6�2��siupdl�]�o�vr�on��`1L�z�`8\�r���il3$|#l4��ǉ#q54Fy�B�Տg{�`���{wc�mס���wxfer��UYtlk2pp<߿UYconv��si�cnv�Qʯxag8��H�Z�lct`ao��=�p��׭nit0�믁�3������  ��� v	��v	$��alFϑpm�r&�B�eWa ���f�%�������I��߬�u�ͬ�Kam�T�f���c��w��ro�ǁ#�5�����?� sm ��y�a��y넑�� ����`����͐ϑ��p��m�Wa�1�� �A�6�S�e�X��ψ� \Q}�����������ĥ w߉�西߭���߮� #q0��rs�ew��� 1�a��z긱n@�.��۲;�d�������  � Ad�	T$�1 p!� P��e �e �	lf@C�@��s/�  ?�����8� ��������reg�.�C=��o9�9 ~@�����$FEAT_IN�DEX  z ���e�� ILECOMP :���1!�!z$#S�ETUP2 ;�1%;"�  �N f!$#_AP2�BCK 1<1)  �)��/�/G  %�/�/e4  �/�/>%�/$?�/H?�/ U?~??�?1?�?�?g? �?�? O2O�?VO�?zO �OO�O?O�OcO�O
_ �O._�OR_d_�O�__ �_�_M_�_q_oo�_ <o�_`o�_mo�o%o�o Io�o�oo�o8J �on�o��3�W �{�"��F��j� |����/�ď֏e��� ���0���T��x�� ����=�ҟa������ ,���P�b�񟆯��� ��K��o�����:� ɯ^�����#���G� ܿ�}�ϡ�6�H�׿ l�����ϝ���@)t �Px/ 2� *�.VR��߅�*��@߂�F�j�T��P�Crߛ߅�FR6�:����V���z�T  �!���K� ��<q�S�*.Fߢ�"��	�Ӑ���^�����STM ��'����S���iP�endant POanelS���HI����9���U�������GIF0;��������JPG��;��]oR�
AR�GNAME.DTy�>�\"����Rc	PANgEL1Y�%>� ��e�w��2�A/@�//���/�3_/��/��/p/�/?�4 �/I?�7?�/?�?�TPEINS.X3ML�?>:\�?t?��1Custom Toolbar�?�Q�PASSWO�RDg?w�FRS�:\:O�? %P�assword ?Config{OR� �OSO�O�O��_�OB_ T_�Ox__�_�_=_�_ a_�_�_�_,o�_Po�_ Io�oo�o9o�o�ooo �o(:�o^�o� #�G�k�� �6��Z�l����� ��ƏU��y������ D�ӏh���a���-� Q���������@�R� �v����)�;�Я_� �����*���N�ݯr� �����7�̿޿m�� ��&ϵ�ǿ\�뿀�� y϶�E���i���ߟ� 4���X�j��ώ�߲� A�S���w����B� ��f��ߊ��+���O� ��������>����� t����'�����]��� ��(��L��p� �5�Yk � $�Z�~� �C�g�/�2/ �V/���//�/?/ �/�/u/
?�/.?@?�/ d?�/�?�?)?�?M?�? q?�?O�?<O�?5OrO O�O%O�O�O[O�OO _&_�OJ_�On_�O_ �_3_�_W_�_�_�_"o �_FoXo�_|oo�o�o��`�$FILE_�DGBCK 1<����`��� ( �)�
SUMMARY�.DG�oblMD�:�o*n`Di�ag Summa�ry+8j
CONSLOG qn��=qConso?le log�7k�pMEMCHECCK��2��q�Memory D�ata3�;g� {�)�HADOW�(�����C�Sh�adow Cha�nges���c-��)	FTP������=��qmment TBD;��;g0<�)ET?HERNET0�`n��q~���=qEth�ernet �pf�iguratio�n��B`%�DCSV�RF/��'�@�C��%� veri?fy allC��c�1p� �DIF�F8��0�ůD�%=Z�diffǯ{���q�1������J�c X�q�|�	�CHGD�&�8�ͿBD�ܯ�����2Ŀ8����R� `�y���GD�.�@���D�q����FY3��8����Z� hρ���GD$�6�H���D������UPDATES.$�
�ck?FRS:\"�c��>qUpdate?s Listc�`{�PSRBWLD.CM��blN��e���pPS_ROBOWEL\�6o+�=�lo a��o����&���J��� n�����9��Jo ���"��X�| #�G�k�d �0�T���/ �C/U/�y//�/�/ >/�/b/�/�/�/-?�/ Q?�/b?�??�?:?�? �?p?O�?)O;O�?_O �?�OO|O�OHO�OlO �O_�O7_�O[_m_�O �_ _�_�_V_�_z_o �_oEo�_io�_zo�o .o�oRo�o�o�o�o AS�ow�*� �`���+��O� �s������8�͏ߏ n����'��� �]�� �������F�۟j��� ���5�ğY�k����� ���B����x������C�үg�v��$FoILE_N�PR]����Y�������MDO?NLY 1<��U�? 
 ��ۿ (���L��5���Y�� }Ϗ�ϳ�B�����x� ߜ�1�C���g��ϋ� ߘ���P���t�	�� ��?���c�u���(� ����^�������$� M���q� �����6��� Z�����%��I[ ���2����?VISBCK����>ų*.VD�*>� FR:\V�� Visio�n VD fileVd����� ��	/./�R/�v/ �//�/;/�/_/q/? �/*?<?�/`?�/�?? �?�?I?�?m?OO�? 8O�?\O�?�?�O!O�O �O�O�O{O_�O!_F_ �Oj_�O�_�_/_�_S_��_w_�_o~�MR_�GRP 1=���LeC4  B�`	 ��lo~l�i`۬B���D��fn���MT� ��� ����e`i`a �o�khb�h�o�dc�ic.N�d��L_L�N�qH���E��|�i`?�{�OA�	�@���=E�{A+8� 3l}�A��A	d�oA	s��sX��p=�l}F@ �qhq��y�~g�fF6��D�MqD��� BT��@���Ô~pD��6����l���5���5��|��~��� B��yB*��B3SlBY�B�B4SM�~T�8�Bp7�aB��A�]wB�Lll叐�A�����A�܏e�P����t����@��bo=���@�	Ƙ����Ο�� +��O�:�_���p������eBH` ������a?���c���'�d
��Z��WZ�m�/��FX
�A@���@��33@�����\��[���ѿ��@ ��񿋯�*��N�9��r�]ϖρ�<�G��=�<�m]�<�+=~�m�<c^��8e�N7��7ѷ7�x7;��51���	ߤ��?ߪ�d2^`Yb`�b`�B���O�i``Үb`� b`�0�����C�^o�߂o�o�߸o ��o�� ]�(߁�l� ������������#� �G�2�k�V�{����� ����������1  ��-�)�� �����0T ?xc����� ��/')�'/M/_/ q/8��/�//�/�/�/ �/?#?
?G?2?k?V? �?z?�?�?�?�?�?O �?1OOUO@ORO�OvO �O�O�O�O��_��J� ���`_*�_N�_�O �_�_�_�_oo'oMo 8oqo\o�o�o�o�o�o �o�o�o7"[F jh�x�t� �!��E�0�B�{�f� ����Ï���ҏ��� �A�,�e�,/������ ���/�J����=� $�a�H�Z��������� ߯ʯ���9�$�]� H���l�����ɿ��ƿ ���#��O�OV� _z� D_V_��z_�Ϟ_�� �
�C�.�g�Rߋ�v� ���߬�����	���-� �Q�<�N��r��� ������)��M� 8�q�\����������� ������7"[F k�|�|���� ֟3�WBg� t�����/� ///S/>/w/b/�/�/ �/�/�/�/�/??=? (?:?s?:�LϦ?p��? �Ϧ� O��$O��T?]O HOZO�O~O�O�O�O�O �O�O_5_ _Y_D_}_ h_�_�_�_�_�_�_�_ o��@o
�go*owo�o �o�o�o�o�o	�o- *cN�r�� �����)�;�M� ��������ˏݏ ď��%��I�4�F� �j�����ǟ���֟ ��!��E�0�i�T��� x���ï�?�?��O� �?OO�t�>O���� ��ѿ��ο��+�� O�:�s�^σϩϔ��� ������� �9�$�6� o�6o��Zo��R����� �����5� �Y�D�}� h������������ �
�C�U��y����� d�����:����� +Q8u`��� ����;& _Jo����� �//گ4/��x�j/ 4��/X�n/|��/��/ �/!??E?0?B?{?f? �?�?�?�?�?�?�?O OAO,OeOPO�OtO�O �O���O�O_�O+__ O_:___�_p_�_�_�_ �_�_�_o ooKo6o ooZo�oZ��o�o�o�o ��xo
G2kR �������� �1��.�g�R���v� ����ӏ���	��-� �Q�/*/��N/��r/ �/ޟ�/��/)�D�M� 8�q�\����������� �گ���7�"�[�F� k���|�����ٿĿ�� �O�O�O��W�B�{�f� �ϊ��Ϯ�������� �A�,�e�P߉�t߆� �ߪ��ߪo��+�=� a��߅�p���� ������� �9�$�]� H���l����������� ����#G2W}�h�p��$FNO ������
F�0� �  #�1 �D|�� RM_�CHKTYP  �� �q�� ��� ��OM� _MsIN� m�����  X� SS�B_CFG >�� �~�Jl�Aj|�T�P_DEF_OW�  m���I�RCOM� ��$�GENOVRD_�DO����T[HR d�d�o_ENB� ��RAVC_GRP� 1?3� X �e/��/�/�/�/�/ �/�/�/? ?=?$?6? s?Z?�?~?�?�?�?�? �?O'OOKO2OoO�O hO�O�O�O�O�O�O��ROU? E� �q������8�?#�O__K_�m_o_ꐖ  D3A���_E�_q�@A��\Bȡ��R��>Y_�6 SMT<#FC-�Ufoxo�o�HOS�TC,1GY?[��_ 	�h�k��o�f�oyeCUgy�z1�������p	�anonymous�5�G�Y�k�w��o �o�o������ *�<��`�r������� ˏ	�����&�8� �������������ȯ گ���M��4�F�X� j�����ݟ��Ŀֿ� ��I�[�m�ρ�fϵ� �ϜϮ�����}���� �,�O�Pߟ�t߆ߘ� �߼���/�A�C�(� w�L�^�p����ϸ� ���������a�6�H� Z�l�~��������� ��9� 2DV�� z������#�� 
.@�������� �������// g</N/`/r/�/�� ��/�/�/?Qcu ��/[?��?�?�?�? �?)/�?O"O4OFOi? �/�/�O�O�O�O9m�a�ENT 1H[� P!^O_  `_?_._c_&_�_ J_�_n_�_�_�_o�_ )o�_Mooqo4o�oXo jo�o�o�o�o�o7 �om0�T�x �����3��W� �{�>���b���Տ�� �������A��e�(��:���^�����㟦�?QUICC0�̟ޟ?��1@��.�����2��l�~�߯!?ROUTER௼��ί/�!PCJO�G0��!19�2.168.0.�10	��GNAME� !�J!RO�BOT���NS_C�FG 1G�I ��Aut�o-starte�d/4FTP:? �Q?SOBχ?f�xϊ� �Ϯ��?�������+� ߿�P�b�t߆ߘ�6 �����(�J� �1� C�U�g�6ߋ����� ����x�	��-�?�Q� c� ?2?D?������� ��)��M_q ����:��� %t�����m�� ��������!/ 3/E/W/z{//�/�/ �/�/�/6HZ ?n/ S?�w?�?�?�?�?�/ �?�?OO<?=O�?aO sO�O�O�O�/
??.? 0O_d?9_K_]_o_�_ PO�_�_�_�_�O�_�_ #o5oGoYoko�O�O�O �O�_�o&_�o1 Cogy����o T��	��-�|o�o �o�o����o��Ϗ� ���)�;�M�_�q� �������˟ݟ�ÿ�T_ERR I������PDUSI�Z  �^����$�>=�WRD �?޵w��  �guest +�}�������ůׯ���SCD_GROU�P 2J� ��`�1��!��L9_���  ��>!�	 i-	�E���Q�E E�ATSWILIB�k�+��ST �4�@��1���L�FRS:аT�TP_AUTH �1K�<!iPendan�������!KAR�EL:*���	��KC�.�@��V�ISION SE!T���u���!�ϣ� �������	��P�'��9߆�]�o޽�CTR/L L��؃��
��FFF�9E3��u���D�EFAULT���FANUC W�eb Server��
��e�w���j��|�������WR�_CONFIG �MY�X�����IDL_CP�U_PC���B��x�6��BH�M�IN'��;�GNR_IO�K���"���NPT_SIM_�DOl�v�TPM�ODNTOLl� >��_PRTY��6���OLNK 1N�ذ�� 2D�Vh��MASTE�k�s�w�OñO_gCFG��	UO��|��CYCLE����_ASG 19O��ձ
 j+ =Oas��������//r�N�UMJ� �J�� I�PCH�x��RTRY_CN�n� ���SCRN_UP)DJ����$� �� ƣP�A��/����$J23_DS/P_EN~��p�~� OBPROC�#ܰ��	JOG�1Q�� @��d8��?� +S? /?>)3POSRE?y��KANJI_� K�l��3��#R����x�5�?�5CL_LF��;"^/�0EYLOGWGIN� q��K1�$��$LANG?UAGE X�6��� vA�LG��"S�߀�����xR��i��@<𬄐�'0u8������MC:\RSCH�\00\��S@N_DISP T��t�w�K�I��LOC���-�DzU�AzCO�GBOOK U 	L0��d���d�d��PXY�_�_�_�_�_� nmh%i��	�kU�Yr�UhozohS_BUFF 1V��|o2s��o�R�� �oq��o�o#,Y Pb������ ����(�U��D/0�DCS Xu] =���"lao�����ˏݏ�3n�IO ;1Y	 �/,����,�<�N�`�t��� ������̟ޟ��� &�8�L�\�n�������ж�ȯܯ�Ee�TM  [d�(�:� L�^�p���������ʿ ܿ� ��$�6�H�Z��l�~ϐϢύd�SE�V� ]�TYP�$���)߄m�1�RSK�!O�c�"FLg 1Z�� ��� �߯���������	�:�STP5@���A]NGNAM�$�E��nk�UPS PGI|%��1�%x�_LOA�D0G %Z%�TEQѼ��MA?XUALRM;'�@I(��~���#� V�#a��CQ[x�8��n���"�1060\	 �F�	�Ϣ������� ������ D'9 ze������ ��R=va �������� *//N/9/r/�/g/�/ �/�/�/�/?�/&?? J?\???�?k?�?�?�? �?�?�?�?"O4OOXO CO|O_OqO�O�O�O�O �O_�O0__T_7_I_ �_u_�_�_�_�_�_o��_,o��D_LDX�DISAc���M�EMO_AP]�E� ?��
  �5i�o�o�o�o�o�o��o��ISC 1]�� �oTd ��\no���� �����I�4�m� �f���$�������� �!��E�ƏT�f�:� ����ß�����z�� ܟA�,�e�w�^���� ��~������ �=� ��L�^�2��������� ߿�r� �Կ9�$�]��o�(t_MSTR �^�͂�SCD 1_xm�W���S��� ����=�(�:�s�^� �߂߻ߦ��������  �9�$�]�H��l�� �����������#�� G�2�W�}�h������� ��������
C. gR�v���� �	�-Q<u `r������ //'/M/8/q/\/�/��/�/�/�/s�MKC_FG `���/~��LTARM_2�a��2 ��#\`Y>G`METsPUT`�"�����NDSP_CMN�Ts506�5�� 	b���>�"1�?�4��5POSCF�7��>PRPM�?�8PSTOL 1c2}{4@p<#�
aA �!aEqOG]OO�O�O �O�O�O_�O�OA_#_ 5_w_Y_k_�_�_�_�_��Q�1SING_C�HK  +O$M/ODAQ73d
?�7�:eDEV 	���	MC:MlHOSIZEs0���eTASK %���%$123456�789 �o�egT�RIG 1e��� l��%��? �  A$�ÜfYP�a,u��cEM_�INF 1f>7� `)�AT&FV0E0�N�})�qE0V�1&A3&B1&�D2&S0&C1�S0=�})ATZ�� �H�E��q9m��xAu���X�������� ���� ��v�)���я��П �������*��N�� ���7�I�[�̯ן�� �9�&���\���� g�����i�ڿ������ ï4��XϏ�iώ�A� ��m�������߿�ѿ B����ϊߜ�O��� ���ߟߩ����>�%� b�t�'ߘ�K�]�o߁� ����(�_�L���p��+����������.ON�ITOR�0G ?�ak   	EOXEC1�#2345�`U789�# ��xxx*x 6xBxNxZxPfxrx22�U2�2�2�2�U2�2�2�2��33�3aR�_GRP_SV �1g�y�a(�Q>`�^�?������ƾee@?�?<I@��Hm�a�_Di�n�!PL_NAME !�5�
 �!Def�ault Per�sonality� (from FwD) �$RR2�� 1h)deX)�dh�
!�1X d �/d/v/�/�/�/�/�/ �/�/??*?<?N?`?�r?�?�?�?�?�?�82 S/�?O O2ODOVOhOzO�O�Ob<�?�O�O �O�O_"_4_F_X_j_�|_�_LhR� 1m�)9`\b0 ��_pb�Q @D7�  �Q?��S�Q�?`�QaAIڏEz  a@og;��	l�R	 0`4b@4c.a�P�Jd�Jd�Ki��K�J����J��J�4�J~��jEa�o�-a�@��o�l[`@��z�b�f�@��S��a�Q�o�c��=�N��
������T;f���`��l[`�*  �p  �$pU> p�$p��o?p?�����O����o�Bn�tr�Q�skse�}�l}�p�  �p�u`j  #p���vks�� 	�'� � ��I� �  {���}:�È6�?È=���N��b@^�d��n�Q��D�{�R�x���nN. ��  '���a�`�@a�@�t��@p@p@C�pC0�f0�+pB�/pC3}�P��@%�Eab�o�o$|m����gA%���. ����z�`�P���QD e���˟��(��m��� �t �O� ru �4 �R�<c��s� :�u�a��P�` �?�f�fb�!�����7� ��گ쬛af�F�>搠���iP�P�;�e�S�Ea4f�u��>LX��s�b<	��I<g�<#��
<2��<D��<��
vo��¯��S��S.���?f7ff?u�?&찗d�@T���?��`?Uȩ?X����Z���T:z�T B��Wa�з*dů�ρ� �ϥ��������&�8�0#�\�h�+�F. K� ��G߼�3���Wɯ�����G�@ G�� ��X�C�|�g�y�� ��������jZ���� ��Q����ߙ����� 3�������/A���t_�����������b���@+Fp�IP��t��%���[`B��0����<ze�xcb!@I�
��M`B@��@�`�9@y��?��h� �@��3�[N��N��N�E��<��/:/L �>���ڟ�A�p�C�F@�S�b/�DpX������@�t��%�h���`/qG���GknF&��FצpE,8{��/ F�ZG����F�nE�DE,ڏ�/�� ���G���F7��F��ED��.��C?.?g? R?d?�?�?�?�?�?�? 	O�?O?O*OcONO�O rO�O�O�O�O�O_�O )__M_8_q_\_�_�_ �_�_�_�_�_o�_7o "o4omoXo�o|o�o�o �o�o�o�o3W B{f����� ����A�,�Q�w� b����������Ώ� ��=�(�a�L���p������(r!3�ji̹�r���ꕢ�3�㱐ڟ�y�4 �����y��P�82�D�&�jb^�p��1w����� ����ʯ���ܯ� �Js�P^�PD�c�`� m���y�\������Ӱ�¿Կ�����.� G����}ϳϡ��� 홍�U�_�J���$�y.�@�v�d�z߈ߚ� x�4�������� ��D�.�2� �$[�G�[�^�B���B��CH� ^���� u�����������p�h�M�_�q�������*���^�^�Y�rm�2��
 �� ��#5GYk} ������h*��� ��>�x}���$MSKCFM�AP  ��� ����m��N"ONREL  6�9_�"EXCFENBkq
7]�FNC��}JOGOVLI�Mkduyd"K�EYk�"R�UN��"S?FSPDTYU��<v_SIGNk}�T1MOT�z�"_CE_GRP� 1n��9\ ���/���/�/4��/? �/2?�/'?h??�?C? �?�?y?�?�?�?O�? @ORO	OvO-OoO�OcO �O�O�O_�O*_<_#_�`_-�"TCOM_�CFG 1o/����_�_�_
|Q_A�RC_�6��U?AP_CPL�_��NOCHECK {?/ 5� ;h9oKo]ooo�o�o�o �o�o�o�o�o#5�GTNO_WAI�T_LF'5y"NT��Qp/���q_7ERR�!2q/_�� R_���"��:�L�dT_M�O�sr�}, ��JP_��_�PARAuM�rs/���`���MW��� =e��345678901.�@�R�)�q���_� ����˟����ݛLW��3�E�؏i�cU�M_RSPACE�,�������$OD�RDSP�SI&�O�FFSET_CAsRToݨDIS��ݢPEN_FIL�E�I!�Q�v�POPTION_IO����PWORK 5t�'� T�|��
� ^�F� �p
���Z���	 �m����A�
��i�_DS�BL  ��v����ޡRIENTkTOj�C����8�ῠUT_SIM_DJ�6	���VàLCT u��}\��Q��W�_P�EXE���RAT����� ���UP� ve������`�����*�8��$���2�#h)deX)�dh�O�X dY�ߑߣߵ����� �����!�3�E�W�i� {������������2n��)�;�M�_�q� ��������<��� ��+=Oas@���X��� O���1m(���(��.�g��"0 �дu�  @D7�  �?���?рH�D4  �EzZ3;�	�l	 0DӀS@SM� �i��i �H)!H�,�H8�H�m�G�	{Gǎ8��6�MV���� �C�)����)����Ճ�*�  �p  �
 > � ,�//�)/ B,�Btr߰«�H�¼�/���/�"`�# �,0 �� _�  � ߽poj  B ��&�X�?MU	'� �� 12I� ��  ���-=����U?g;/�@}?�0~.ѱ�?;Ѳ����H[N5��? � 'M�D�> C)�f)�J BN +��=x%O7O�R�@D1~�oo$�����JWA�D0�J5�4�:  �1�E&?�O�O#_�_G_2]�� ��t O� �ru �4 ���R�Uɳ� :��%Ёр� �?�ff��@[�_�_BV_{�o~��18р�"o0j>�P�Q6YP�рZo�WrAdS�%��>Lw0�#�<	��I<g�<#��
<2��<D��<�׍�l��_�ѳMb�@?offf?�0?&p�:T@T�q?��`?Uȩ?X�-q�iyBq5Y a��gI�_� �����!��E� W�B�{���d�����Տ�LnpΏ/�ʈG�@ G��U�ȏy� d�������ӟ����� ��yB=� ��?p�� �/򏸯�߯R��� '�9��oN�`�����~�P����ۿƿ�B�� �D�e�ֿ;�ҿ_�J�?��h�oϨϓ�J���D4��b!�_@ ���� ߧ��Ŀ�����%�@I�)�M`�B@��@`��9@y��?��h	� �@�3��[N��N�N��E��<�/�Y�kЖ>��ڟ��A�p�C��F@�S���pX������@��t��%�h���߉!G��G�knF&�F׿�pE,8{�� �F�ZG����F�nE��DE,ڏ������G��F7���F��ED��Mf��b�M��q�� ����������(�� 8�^�I���m������� ��������$H3 lW�{���� ��2VAS �w������ /.//R/=/v/a/�/ �/�/�/�/�/�/?? <?'?`?K?p?�?�?�? �?�?�?O�?&OO#O \OGO�OkO�O�O�O�N=(]�3�ji�O�a���	U�E3Ա�x�O_<q4 ��%_<7_<q�P�Q_c_�ERjb}_�_1w?������]�Y��_�_o�_1ol��P�bPcn~���o�O@�o{_�o�oY�`��o �o,/;M#�f 0o�����Y�e@t�~�i#�1�C�yM� _�����������{bS� Ԏ��	�?�-�c�Mj�2���$�VG�Dz}�B����B��CH�}�9�֟��� ��0�B���wl�@~�������Ư�T�E��\��qQ��U
 ί�0�B� T�f�x���������ҿ����χ��� ���]{x}��$P�ARAM_MEN�U ?Յ��  �DEFPULSE��	WAITT�MOUTl�RC�V� SHE�LL_WRK.$�CUR_STYLvj���OPT��N��PTB����C��R_DECSNw� Te'�!�3�E�n�i�{� �߶߱������������F�A�USE_P�ROG %P�%�B��V�CCR���UeXÚ�_HOST7 !P�!����Tt`����������4���_TIME��� �T�  A�GDEBUG��P�V��GINP_FLM3SK]���TR����WPGA�� |�[����CH����TYPEM�Y�A�;�Q zu������ 
)RM_q �������/ */%/7/I/r/m//�/��/�/�/�/?��WO�RD ?	��	�RS��CPNeS�E��>2JO��ξBTE���TR?ACECTL�PՅ�Z� {`�/ a`{`�>�q6DT QxՅ��0�0D��Sc7{a�0����2���?�?�2��4D�2#A�O.O@ORFcA�bBU`D	`D
`D`DU`D`D`D`DU`D`D`DObOtO�F A�5P�2 Q0TOBPRPBP�BP0T�BP�BP�BP�A,_>Z�_=_ O_a_s^$_�_�_
b�� "o4d�_�_�_�O�O_P_a�1	ad�TUVd^dfdnb�Wr�k}�o�o��j;qwc�TvT ~T5OcM_q�� ���v,>�
�t �@�R�d�v������� ��+������ˏ�� u������ԟ����9�*�<�N�`� r���������̯ޯ� ��&�8�J�\�n��� ������ȿڿ���� "�4�F�X�j�|ώϠ� ������������0� B�T�f�xߊߜ߮��� ��������,�>�P� b�t��������� ����(�:�L�^�p� ��������������  $6�Fl~� ������  2DVhz��� ����
//./@/ R/d/v/�/�/�/�/�/ �/�/??*?<?N?`? r?�?�?�?�?�?�?�? OO&O8OJO\OnO�O �O�O�O�O�O�O�O_ "_4_F_X_j_|_�_�_ �_�_�_�_�_oo0o BoTofoxoN�o�o�o �o�o�o,>P bt������ ���(�:�L�^�p� ��������ʏ܏� � �$�6�H�Z�l�~��� ����Ɵ؟���� � 2�D�V�h�z������� ¯ԯ���
��.�@� R�d�v���������п �����*�<�N�`��rτϖϨϺ����$�PGTRACEL�EN  ��  ��������_UP y/�����������_CFG7 z�����e��<��� <��Z�l�<�$�DEFS_PD {/��a������IN'�T�RL |/�S�8�Lԃ�IPE_CO�NFI+�}����<�x�L�ID(�~/��G�RP 1���������@�
=��[���A?C��C
�XC)���B��r�������dL�z������� 	 r�N������ ´����B������������A���> �6>7��D_������� ='�=)��� ������	B-���Q�M���  #Dz����
� �&L7p[� �����/�6/�!/Z/��
V7.10beta1<�}� B=q�"�`ff@��">�����!=���ޏ!A>ff�!@ֻff�"�\)�"D���?�  �!@��!� �!Ap�#W���h/??*?<?K;�w����O/�?K/�? �?�?�?O�?O>O)O bOMO�OqO�O�O�O�O �O_�O(__L_7_p_ [_m_�_�_�_��_ o �_$oo!oZoEo~oio �o�o�o�o�o�o�o �DQy{/�#F@ {yw}�y{ջy�- ������/�Z?l? ~?w���t�����я�� �������O�:�s� ^���������ߟ�ܟ � �9�$�]�H���l� ~����_ۯ����� 5� �2�k�V���z��� ��׿¿�����1�\ n�j�|϶���� ���	�4�F�X�j�c� χߙ߄߽ߨ����� ���)��&�_�J�� n����������� %��I�4�m�X����� ί����������! E0B{f��� ���H�Zό� Vh�ϴϊ���� � �2�D�V�O/�s/ ^/�/�/�/�/�/�/�/ ? ?9?$?6?o?Z?�? ~?�?�?�?�?�?O�? 5O OYODO}O�O���O �OtO�O�O_�O1__ U_@_R_�_v_�_�_�_ �_�_"4FxBo| ����o��o�o/ /0/B/;�__J� n������� %��I�4�F��j��� ��Ǐ���֏�!�� E�0�i��O^���N�ß ՟�������A�,� e�P�b���������� o o2oTo.�hozo�o �����o��Ϳ�o
 گ'�֯K�6�o�Zϓ� ~Ϸ��ϴ�������� 5� �Y�D�Vߏ�z߳� �����������1�� Uy��:����� ����	���-��Q�<� u�`�r���������� �T�f�x�n� ���������� �7"[Fj� ������!// E/0/i/T/f/�/�/�/ �/�/�/?�//?A?l� e?w?&?�?�?�?�?�? �?�?OO=O(OaOLO �OpO�O�O����*�O�_@RdZ_l_���$PLID_KNOW_M  �?��A�T�SV ��.�P�[?�_ �_o�O&oo#o\o�B���SM_GRP S1��Z� dI`�?oo$Cf�d�����D� �TPbj�oLk�f�o"~ �U�o>n2T �~�����7� 4���p�D���R��� ʏ����������6�
��T��*������QMR��c��mT�EGQK? GR��(�#���[� �/�A�S��������� ���$����W��+� =�O������������� ���S�Ͻ�ST^�a1 1�������P0� @� ���E�ϲ�������� �M�0�B�T�fߧߊ� ������������7��(,�m��2�����A'�<��z�3��������4����������5)�;�M�_���6 x���������7����������8(:L~��MAD  ����� ��PARN_UM  ��Ko\���SCH�
 ��
��S+UP�D��xaq{��_CMP_�`� <Pz �'�U�ER_C;HK����Z����RS���_�Q_#MO� �%_���_RES_G����� ��v/{/�/�/ �/�/�/�/�/*??N?�A?r?e?w?J'��W, g/�?L%��?�?�?N# (��?OON#w�4OSO XON#��sO�O�ON#  �O�O�ON#d �O__N"V 1��Uua��@cX��Pp�P$�@cW،P��P@�@cV��P�"T?HR_INR����pbA%d�VMASS6�_ Z�WMN�_�S�MON_QUEU�E ��e��`Ȫ�`�N�U�N8�V�2`END4a6/�NiEXE]oNeWB�E\`>o/cOPTI�O;g?+2`PROG�RAM %j%�1`O_�0bTAS�K_I��nOCFG �o�9p�DATAɓ�B{@ev2w���� ��z��+�=�O���s���������nzIN+FOɓ��}�!dr� �!�3�E�W�i�{��� ����ß՟������/�A�S�e�w�҇ބ�Ɔ| �98q�DI�T �Bׯj~W�ERFL~hwS~�RGADJ �ƪ/A�  ,�?E�8���Q�IORITY��W���MPDSQP�a�j�U�WvTv�OG��_TG����Rj��TOE�P1��ƫ (!A�F�PE5 ���!�tcp��%�!�ud�?�!i�cm<�Q_��XY_�<q�Ƭ�Oq)�� *������Op������������<� #�5�r�Yߖ�}ߺ��ߠ�������&�*�P�ORT�a�Op�A%�_CART�REP~`Ʈ��SK�STA�X!*SSA�V`�ƪ	25?00H809u�T�毙䕣�ƫ�����`X#�$�6�m�/URGEU`B��A)WFP�DO�V�2��W�q�?Q�WRU�P_DELAY ��Ưe�R_HO�T�hwR%z����R_NORMAL�nx��6SEMI�:y�QSKIPڕ��X%�x 	������� �X%-;%[m E������� !//E/W/i///y/�/ �/�/�/�/�/?�/? A?S?e?+?�?w?�?�? �?�?�?O�?+O=OOO�1U�$RBTIF|��NaRCVTM��v���m@DCR�햜�A@&�HB�-�AȤ��@=ʄ@��߰)܀���d{sJ/ž
�n�Ꮹ�|�_ �<	�I<g��<#�
<2���<D��<��
+__{_�_)`���_ �_�_�_�_ oo$o6o HoZolo~oi_�o�o�o �o�o�o�o DV �_z������ �
��.�@�R�=v� a�����������׏ �*�mN�`�r����� ����̟ޟ����� 8�J�5�n�Y���}��� ȯ�����A�"�4�F� X�j�|�������Ŀֿ �ӯ���0�B�-�f� Qϊ�m��������� ��,�>�P�b�t߆� �ߪ߼ߧ�������� (�:�%�^�A����� �������� ��$�6� H�Z�l�~���{���� �������� 2V h������� �
.@R=O �s�����/ �*/</`/r/�/�/ �/�/�/�/�/??&?�28�AGN_ATC� 1��K �AT&FV0E�02;ATDP�/6/9/2/9�p8ATA2>,�AT%G1%�B960k9+�++�?,�1H�?,��AIO_TYPE'  EC/4?�REFPOS1 �1� K x�O[H/O/�O�M NO`O�O�O�O_�OC_��Og__d_�_+K2 1� KLON_�_o��_*o�_5A3 1� �_�_�_ o�o�o�o@oS4 1�Woio{o�o3W�oS5 1��o�oJ��|�jS6 1������]�H����S7 1��(�:�t���ݏ���S8 1�����Ϗ	���r����)�SMASK 1� O  
���ɗ'XNO�?���1.��8�1AMOTE  ��.DN�_CFG ��U���5�0BPL_RANGQ�K!Y��POWER ��Q5 a�SM_D�RYPRG %��%R���ȥTAR�T ����UME_PROׯ�d��.D_EXEC_E�NB  �5]�GSPD=����Y3��gTDB����RMÿ.��MT_ѐT��S��D0OBOT_N�AME ��S�;9OB_ORD_NUM ?���AH80�0I$�	��se	�\������ ��e��	@��}�D|��D0PC_TIMEOUT��{ xD0S232n��1�Q; L�TEACH PE�NDAN��j�5���=Q�x0Mai�ntenance ConsK"-���"+�t4KCL/)C�}�6��|�� No Us�e�=[߹�F���NPqO�ќ�5�_����CH_L@���U���	J��MAVAIL`���+���]�I�SPACE�1 2�=L �����p��扢�J@����8�? ��� ���V�w�N� �������������� 4�&G
l�}d	Q5 U1���������` 4&G
l}d�#��2������ ��2A/b/%/w/�//�/�3��� �	/�/-/O/^??B? �?�?�?�?�4�/�/ ??&?�?J?l?{O�O@_O�O�O�O�O�5�? OO1OCO�OgO�O�_��_|_�_�_�_o�6 _*_<_N_`_o�_�_ �o�o�o�o�o!�75oGoYoko}o+�o �o����)��>��8Rdv��H� ����ӏ%�F�-��[��G ��� R�;�
�� ����ԟ���
�� .�@����c���p���8�¯=�dؠ��ϟ�� �!�3�E�W�i�_�q� �����x��կ�� '�9�K�]�oρ�w��� ����Ͽѿ����5� G�Y�k�}ߏߡߗ���p������� `S� @��8堯F�"�*ل������ �������,���� V�h�2�<�N������� ������.L4 v�R\n�����
f�7�_MO�DE  ��MS ���&����AÏb��*	��&/�$CWORK_{AD]	)`\�!/R  ���t �+/^ _INTVA�L]���hR_O�PTION�& �h�$SCAN�_TIM\.�h��!R �(�3�0(�L8������!��3��1��/@>.?����S22�41�9dD�4�1"3��@��@�?�?�?���IP���@���JO8\OnOE@D���O �O�O�O�O�O__(_�:_L_O���4�X_�_�_��8�1���;�o�� 1��p�c]�t��D�i�1��  � lS2��15 17oIo [omoo�o�o�o�o�o �o�o!3EWi {����wc�� �	��-�?�Q�c�u� ��������Ϗ��� �)�;�M�_���`[ ����ğ֟����� 0�B�T�f�x������� ��ү�����$�7�  0��� om�� ������ǿٿ���� !�3�E�W�i�{ύϟ� ��������v���/� A�S�e�w߉ߛ߭߿� ��������+�=�O� a�s�����ߖ��� �� ��$�6�H�Z�l� ~���������������� 2DVP�\�  �A������ �%7I[m �������/ �/C(/N/ `/r/�/�/�/�/�/�/�/?F;/?B?F;�x1 ;?w=�	123456�78{��
l�@�P�?�?�?�?�?O9/2ODOVO hOzO�O�O�O�O�O�O -/
__._@_R_d_v_ �_�_�_�_�_�O�_o o*o<oNo`oro�o�o �o�o�_�o�o& 8J\n���o� �����"�4�F� X�j�|������ď֏ �����0�B�T�f� ����������ҟ��� ��,�>�m�b�t��� ������ί����(��6yI�[�@�`����������Cz � Bp*   ���254F��$S�CR_GRP 1��(�e@(�l߀�0@� `1 �[1s	 )�3�C�<�t� vrY�8P�}�kϤ�n���95C�����-u��ȡ����LR Mate 200iC �1�90�1Շ0LR2C �3�=OÆ�ED�
f؜1u�2�@U7��`1��v��@�u���	t��������4�$�^0�2��� _2T�gϡϊ��o�F� D�f?��s�����￶}ht ,Z�mo| -ON�B�˰�P�N��g�N�Aܰv�  @�DЎ�N�@����  ?� ��J�H˰��y��N�F@ F�` ������A,Q wb���n�N���������B� �_J�n�� ���/�%//I/ ��E+:3��6?|?�5�ա
�/�/�#��@=���"�/pǢ� 3Bm�07�590@7����EL_DEFAULT  I���� �^1MIPOWERFL  V�v5]2ރ0WFDOk6 �v5 �ERVENT? 1���O�t3�C�L!DUM�_EIP?�8�j�!AF_INExj0O�$!FT�?�=NOaO!Q�O ��PO�O!RP?C_MAIN�O�Hq��O�O�CVIS�O�I��OE_!TP&8PPU<_�9d4_�_�!
PMON_POROXY�_�6e�_��_XR�_�=f�_)o!�RDM_SRV�*o�9gouo!R�R8�o�4hdo�o!
��@M�_�<i�o!RLSYNC�4y8�oY!R3OS�?�|�4H� tO�8c����� ;��_�&���J���n� �����ȏڏ7�I���m�4���X����7I�CE_KL ?%��; (%SVCPRG1���안�!��3*�/��4�R�W��5z���6�����7ʯϯ�C�$�5�9��o G����o������ D����l��񑔯� 񑼯7���_��� ���4����]���� �������'��տO� ���w��%ϟ��M� ���u�������� ��?�A��Ͽ�ђ�؟ ꐊ���ɱ������� �?�*�c�N������� ����������) ;_J�n��� ���%I4 mX�|���� �/�3//W/i/T/ �/x/�/�/�/�/�/�/�?/??S?Ś_DE�V �9��MC:[8�i.m4OUT_Rf1~6~i8REC 1����f0�0 �1 	 �2�?�1���3O�MO@O+OdO��
 ��Z���6 �s  UEBf0KX�q�0�0�f0ʬ��2�3f0nf0�@ ���-�X�O�2E0��0'qE0_�O_�5 "_�C&_L_:_p_^_�_ �_�_�_�_�_�_o o "oHo6oloNo`o�o�o �o�o�o�o D 2TVh���� ����
�@�.�P� v�X�������Џ��� ��*��N�<�r�`� ������̟��ܟޟ� &��J�8�n���b��� ��ȯ��دگ�"��3 ~A�(��P���t��� ��ο�¿��(�� 8�:�Lς�dϒϸϦ� ���� ���$�6��Z� H�~�lߎߴߢ��ߺ� �����2� �V�D�z� ��n���������
� ��.�@�"�d�R���v� ������������ <*`N��x� ����8 HJ\�������G�5V 1��< �P_�1��FO�2�  j�0eXF>a?_TYPE�?k2�HELL_CFG� �z:f2/ ��B�/�/ %RSR�/�/�/?
?C? .?g?R?�?v?�?�?�?��?�?	O�?-O?O/�  �!�@oO�OP�O�C�I�AP�OL�B�@�WgB2P�d�O�O�&HK 1��+ �OE_@_ R_d_�_�_�_�_�_�_ �_�_oo*o<oeo`o�ro�oa&�#OMM ���/�o�"FTOV_ENBr$!}*�OW_REG_U�I�oe"IMWAI�T�b�I${OUTrv$&yTIMuw��`VAL5>'s_UNIT�c�v�})MON_ALI�AS ?e�i ( he!� �� $�6�Q&�c�u����� D���Ϗ�����)� ;�M�_�q�������� ˟ݟ����%�7�� H�m������N�ǯٯ ������3�E�W�i� {�&�����ÿտ習� ��/�A��e�wω� �ϭ�X��������� ��=�O�a�s߅�0ߩ� �����ߊ����'�9� K���o�����b� �������#���G�Y� k�}���:��������� ��1CU y ����l��	 -�Qcu�2 ������/)/ ;/M/_/
/�/�/�/�/ �/v/�/??%?7?�/ [?m??�?<?�?�?�? �?�?�?!O3OEOWOiO O�O�O�O�O�O�O�O __/_�O@_e_w_�_ �_F_�_�_�_�_o�_ +o=oOoaosoo�o�o �o�o�o�o'9 �o]o���P�������s�$S�MON_DEFP�RO ����:� �*SYSTEM*  �l�*��RECALL ?�}:� ( �}�5xcopy f�r:\*.* v�irt:\tmp�back��=>l�aptop-u9�nqdgeh:5�928 ��3 723 5�͏ߏ�s}6z�a���������B�T��:{�s:o�rderfil.dat������ӟ��}1{�mdb: �������=�O�a�� y�������ү��� ����-�>�P�b�u��� �����ο����� )���L�^�q����� 9���������%��� H�Z�m����5��� �������!ϳ�D�V� i�{�ߟ�1�����g� �ϊ��/�@�R�d�w� ���-�������ߐ� ��+�<N`s��� ��;�����'� �J\o���
��7 �������#�F/ X/k}�3/�/�/ ���/�/�/B?T?�/ y�///�?�?�?� �?/�?>OPObOu/? O�/�O�O�O�/�O�O )?�OL_^_q?�?O�? 9_�_�_�?O�_%O�_ HoZomOO_�O5o�o �o�O�O�o!_�oDV i_{_�_1��g �_�o�@�R�d�wo 
��o��Џ��o�����+<�N�`�ss
x�yzrate 61 ��)�;�̟ޟ�qu!z���39020 ����?�Q�c�vp�tpdisc 0���,���ϯ��trtpconn 0 ��������J�\�ow;z����6�ǿٿlz2�������>�P�b�op�$SN�PX_ASG 1߶������� P�'�%R[1]@g1.1f�ly?�os%���Ͽ� �����6� �@�l�Oߐ�s߅��� �������� ���V� 9�`��o������ �������@�#�5�v� Y������������� ��<`CU� y������& 	0\?�cu� ����/�/F/ )/P/|/_/�/�/�/�/ �/�/?�/0??%?f? I?p?�??�?�?�?�? �? O,OOPO3OEO�O iO�O�O�O�O�O�O_ �O _L_/_p_S_e_�_ �_�_�_�_ o�_�_6o o@oloOo�oso�o�o �o�o�o�o V 9`�o���� ����@�#�5�v� Y�������Џ��ŏ� ��<��`�C�U��� y���̟���ӟ�&� 	�0�\�?���c�u��� �����ϯ���F��)�P�|�_�x�PAR�AM ������ �	���P���p�OFT�_KB_CFG � ����״PIN_SIM  �ˁ̶�/�A�ϰx�R�VQSTP_DS�B�̲}Ϻ���S�R �	�� &� TEST V����ԶTOP�_ON_ERR � �����PT�N 	���A��RINGo_PRM�� ���VDT_GRP �1�����  	 з��b�t߆ߘߪ߼� �������+�(�:�L� ^�p��������� �� ��$�6�H�Z�l� ~���������������  2DV}z� ������
 C@Rdv��� ���	///*/</ N/`/r/�/�/�/�/�/ �/�/??&?8?J?\? n?�?�?�?�?�?�?�? �?O"O4O[OXOjO|O �O�O�O�O�O�O�O!_ _0_B_T_f_x_�_�_ �_�_�_�_�_oo,o >oPoboto�o�o�o�o �o�o�o(:L sp�������� ��9�6�׳VP�RG_COUNT������d�EN�B/�_�M��鴖�_�UPD 1�	�8  
M������ �-�(�:�L�u�p��� ������ʟܟ� �� $�M�H�Z�l������� ��ݯد���%� �2� D�m�h�z�������¿ Կ����
��E�@�R� dύψϚϬ������� ����*�<�e�`�r� �߭ߨߺ�������\�YSDEBUGn��Ӏ���d��"�SP�_PASSn�B�?4�LOG �V΅�������
�  �����
�MC:\`��a�_MPCf�΅����ҁ���� ҁ��SA/V �i��������SV�T�EM_TIME �1�΋ (u���q�������T1S�VGUNSɀo�'������ASK_?OPTIONn�΅�������BCCFG �΋O���I�2��`;A�I�r ]o������ �8J5nY� }�����/� 4//X/C/|/g/�/�/���,�/�/ ??�/ �/H?3?l?W?�?��? ��0�?�?�?O�?&O OJO8OZO\OnO�O�O �O�O�O�O_�O _F_ 4_j_X_�_|_�_�_�_ �_�_o�X�  o2oPo boto�_�o�o�o�o�o �o�o:(^L �p����� � �$��H�6�X�~�l� ����Ə���؏���� �D�2�h�o������ ԟR�����.�� R�d�v�D��������� �Я����<�*�`� N���r�������޿̿ ��&��J�8�Z�\� nϤϒ���~������ "�4߲�X�F�hߎ�|� �����ߤ������� B�0�R�T�f����� ����������>�,� b�P���t��������� ����(��@Rp ������� $6ZH~l ������� / /D/2/h/V/x/�/�/ �/�/�/�/
?�/?? .?d?R?�?>�?�?�? �?�?r?OO(ONO<O rO�O�OdO�O�O�O�O _�O__&_\_J_�_ n_�_�_�_�_�_�_�_ "ooFo4ojoXozo|o �o�o�o�o�? 0 BT�oxf��� ������>�,� b�P�r�t��������� Ώ��(��8�^�L� ��p�����ʟ��ڟܟ �$��H��o`�r��� ����2�دƯ�����2��P��$TBC�SG_GRP 2���� � �P� 
 ?�  {���w��� ��տ��ѿ���/�A��T�[��b�d0� �p�?P�	 H;BHA�L�͌�@�B   C���϶˘���ϟ�D����AQ���x���A��T$��9��6ff��f�@2P�C�ώ�@�f߬��C��ߐ߮ߴޥ� ��%��%�D�W�"�4��j�|�������?�Y�����	�V3.00s�	�lr2c��	*�2�*�O�A� ��ѳ3e3P�d��� x�J�y�  �������T�JCFG Ė�l� o������������=K
%�Kq\ ������� �7"[Fj� ������!// E/0/i/T/f/�/�/�/ �/�/�/s���??(? �/[?F?k?�?|?�?�? �?�?�?O!O3O�?WO BO{OfO�O�OP�<��O ��O�O�O0__T_B_ x_f_�_�_�_�_�_�_ �_oo>o,oNoPobo �o�o�o�o�o�o�o :(^L���� ��h� ��$�� H�6�l�Z�|�����Ə ��֏؏� ��D�V� h�z�4�������ҟ ԟ��
�@�.�d�R� ��v��������Я� ��*��:�<�N���r� ����̿���޿ �&� �>�P�b�ϒπϢ� �϶��������4�F� X�j�(ߎ�|߲ߠ��� ��������B�0�f� T��x�������� ���,��P�>�t�b� �������������� &(:p^�� ��t�����6 $ZH~l��� ����/2/ /V/ D/z/�/�/�/j/�/�/ �/�/?.??R?@?v? d?�?�?�?�?�?�?�? OO<O*O`ONOpO�O �O�O�O�O�O_�O_ _&_\_�t_�_�_B_ �_�_�_�_�_"ooFo 4ojo|o�o�o^o�o�o �o�o�o0B�o xf������ ���>�,�b�P��� t���������Ώ�� (��L�:�\���p��� ��ʟ��� ��_�*� �_�l�Z���~����� į�د� �2��� h�V���z���¿Կ� ��
�����.�d�R� ��vϬϚ��Ͼ���� ��*��N�<�r�`߂� �ߖ��ߺ������� 8�&�H�n�\���>� ����x������4�"� X�F�|�j��������� ������
Tf x�D����� �P>tb �������/ /:/(/^/L/n/p/�/ �/�/�/�/ ?�/$?6? ��N?`?r??�?�?�? �?�?�?�? OODOVO hOzO8O�O�O�O�O�O��N  PS �V$_R�$TB�JOP_GRP �2��E�?  ?�W<R�CS�J\��@�0WP�R@T�P ט ��T�T ��Q[R	 �BL�  �UCр D�*W[Q�_�_?ff�fe:lB ��P�ff@`�?33D  $a�U 3o>g�_�_po�l�P�e�9<�bbY���?٪``$o�oUAm��gD�`$�co�Quz9�P��Aa�P@a����C�Z`Ep�o]A63ffpu`aD/�U�h�͔r��~�a�R@ieAq�`�q��@9q�|�d&`%���c�333D�\P8���?�`?L�pAp[QB�b�k�}� ��z>�� >�ffԁL���T�f��fo � �Nw@�*�8�f���r� ,���П��ȟ��'�� ��F�`�J�X�����S�C�Vء��	�V3.00�Sl7r2c�T*��T�Q�� E����E�A E���E��3E��iNE�!hE��فEۑ�E��I�E��E����E�rF��F�F�M(F�5F�BFaOF��\F"f,�z�  E�@ E��� E�� E��  E����� �E����� E�ꆰԎ�ᆰ� �F   F� �F$ Fj` �F�@ F�P �F�` 9�IR/9�o���L�Q_ ��V���LQ�8TESTP�ARS�XUP9SH�Rk�ABLE 1%�J[4�SV�+�Q �0�V�V�VȨWQV�	V�
V��Vȥ�QV�V�8V�뱅�RDI��TQ�϶���������f�On߀ۊߜ߮�������Sl�RS 0ړ�� �����������#�5� G�Y�k�}��������� ����/]k�o��*	� %�7�I�����+�=��O؆�NUM  ��ETQ�P�P �밆�_CF�G ����Q@�<PIMEBF_T�Tq��RS~�;VE�R�<Q;R {1�J[
 8��RP� �@5  ������/ /&/8/J/\/n/�/�/ �/�/�/�/#?�/?Y?@4?F?\?j?|?{_��h@R
<PMI_�CHANG R >�3DBGLVQ`I�R;Q�0ETHE�RAD ?�E
;@�S �?�?TO6V��0ROUTe!�JZ!�D�OwLSN�MASK0HRSAA255.�E��O�O�8TOOLOFS_�DIq��5IOR�QCTRL �s[���n]8]_�_�_ �_�_�_�_�_o"o4o�Fo�
�_Tofo�og�PE_DETAIH�3ZPON_SVO�FF)_�cP_MOON �"P2�i�STRTCHK ��J^mO�bVT?COMPAT�h;C��d�`FPROG %JZ%j�=?~qqISPLAYr���j_INST_M��@ �|�g�tUS8e]orLCK��{QUICKME�0�)�orSCREF�}3Jtps��@or�a�f��2w�_{����ZyISR_GR�P 1�JY ؛ 6���@��;�)�_�M��8 ����Y�������͕ �����/��S�A�w� e�������ѯ��������=�+�M�s�	�12345678h����f�X`�1�Ћ�
 �}ipn�l/۰gen.htm�����0�B��X�Panel� setupF�}�<�ϘϪϼ����� u�k��*�<�N�`� r��ϖ�ߺ������� ��ߝ�J�\�n�� ����I�?������ "�4�F���j������ ��������_�q�0 BTfx��� ����>� bt����3�~�UALRM�pG {?J[
  � */!/R/E/v/i/�/ �/�/�/�/�/�/??�<?�SEV  ��n6�ECF�G ��m�6��A��1   Bȩt
 =?�s3E�?�?�? OO+O=OOOaOsO�Oh�Gz1ʂ��k S(Ο�OH7Isv?}{�`(%0?"_p_I_4_ m_X_�_|_�_�_�_�_��_o�_3o�L� ��M�OAoI_E�HI��p1��i  �( k`��(/�SOFTPART�/GENLINK�?current�=menupage,153,1}o0�o&�'�o�n71�oq���6qy);�eedit�bT��`�	��-�8Je,2�ox������=��oT�148,A2�� ��$�6��)o [�m��������D�ٟ ����!�3�W�i� {�������î�R��a R����%�7�I�L� m��������ǿV�� ���!�3�E�Կ�{� �ϟϱ�����d���� �/�A�S���w߉ߛ� �߿���`�r���+� =�O�a��߅���� ����ʯܯ�'�9�K� ]�o�r���������� ��|�#5GYk }������ �1CUgy ������	/� -/?/Q/c/u/�//�/ �/�/�/�/?���;? M?_?q?�?�?�/�?�? �?�?OO�?7OIO[O mOO�O�O2O�O�O�O �O_!_�OE_W_i_{_ �_�_._�_�_�_�_o o/o�_Soeowo�o�o �o<o�o�o�o+ ?(?as���� �o����'�9�� �o���������ɏX� ����#�5�G�֏k� }�������şT�f��� ��1�C�U��y��� ������ӯb���	���-�?�Q�<��$U�I_PANEDA�TA 1�������  �	�}/fr�h/cgtp/w�holedev.stmc���ӿ���>�)pri��.�Ip}2�V�h�zόϞ��� )���Ͻ����� �0��T�;�xߊ�q߀�ߕ��������Bv�Nq*�=�B�T� f�x�������3��� ����,�>�P���t� [�������������� (L3p�i�� �������� �1C�g�� ������L	/ //?/&/c/u/\/�/ �/�/�/�/�/�/?�/ ;?M?���?�?�?�? �?�?0?Ot%O7OIO [OmOO�O�?�O�O�O �O�O_�O3__W_i_ P_�_t_�_�_�_�_Z? l?o/oAoSoeowo�_ �o�o O�o�o�o +�oO6s�l� ������'�9�  �]�D����_o�oɏ ۏ����#�v�G��o k�}�������ş,�� �����C�U�<�y� `�������ӯ����ޯ �-�����c�u����� ������T���)� ;�M�_�q�ؿ��|Ϲ� �����������7�I� 0�m�Tߑߣߊ���:� L����!�3�E�W�� {�� ϱ��������� �r�/��S�e�L��� p������������ =$a����}��r�����) �*��Vhz� ������� .//R/9/v/�/o/�/ �/�/�/�/?��������$UI_PAN�ELINK 1����  ��  ��}�1234567890_?q?�?�?�?�? �4��]?�?�?OO1O CO�?gOyO�O�O�O�ODYIY0:�M��[0�-/SOFTPA�RT/GENA1?�CONFIG=S�INGLE&PR�IM=mainedit �OI_[_m_�YJ_$_M=wintpe,1@_�_�_�_XK  �_$o6oHo Zolooo�o�o�o�o �o�o�o
2DVh z������ ��.�@�R�d�v���  �����Џ����M� 0,M9P �E=Por?S�,Ico:�{�^����� ��˟ݟ�����7�@�[�m�P������O����BS0ߢ��C�� �/�%�7�I�[�m�`C �������Ϳ߿񿀿 �'�9�K�]�o��L�� �э͙�Q|������� ���!ߨ�;�M�_�q� �ߕߧ�6�������� �%��I�[�m��� ��2����������!� 3���W�i�{������� @�������/�� Sew����.� ��z�!E( W{^����� �/�//A/���͡� ��}����/�/�/�/�/ ?�2?D?V?h?z?�? ?�?�?�?�?�?
OO �ϝϯ�dOvO�O�O�O �OE�O�O__*_<_ N_�Or_�_�_�_�_�_ [_�_oo&o8oJo�_ no�o�o�o�o�o�oio �o"4FX�o| �����e�� �0�B�T�f����/ ���������ُ��� >�P�3�t���i����� Ο��O/�s/(��/L� ^�p����������?ܯ � ��$�6�ůZ�l� ~�������#O5OGO� � �2�D�V�h���� �ϰ�������u�
�� .�@�R�d�v�ߚ߬� �������߃��*�<� N�`�r������� �������&�8�J�\� n�������������� ��m�"4ßXjM �q������ BT7x��� ���A��//,/ >/P/C�t/�/�/�/�/ �/�/o/??(?:?L? ^?Ϳ߿�?�?�?�? �? OO�?6OHOZOlO ~O�OO�O�O�O�O�O _�O2_D_V_h_z_�_ �_-_�_�_�_�_
oo �_@oRodovo�o�o)o �o�o�o�o*�o N`r���� �m��&�8��\� n�Q���u���ȏ��� ���"���?�?�{���$UI_POSTYPE  �5� 	k��{��_QUICKMEN  ���j�����RESTO�RE 1ו5�  � �/
�2�D�h�mc��� ����¯ԯw���
�� .�@��d�v������� W���˿ݿO��*�<� N�`�τϖϨϺ��� �ρ���&�8�J��� W�i�{��϶������� �ߡ�"�4�F�X�j�� ��������ߋ��� �y�+�T�f�x����� ?�����������, >Pbt���� ��(�L ^p���I���� //��SCRE�ܐ?�uw1sc-�u2M$U3M$4M$5M$6M$�7M$8M!��USE�R/ 4/F"T. O#k�sW#�$4�$5�$6ʶ$7�$8�!��ND�O_CFG ض��  ,� ��P�DATE �)��None �V��SEUFRA_ME  
��&�,1RTOL_AB�RT7?��N3ENB�X?I8GRP 1��!��Cz  A��3�1��?�?�?�?��?FO"OG:ېU�x81g;MSK  �{5�Ag;N41%�a��B%��O��VI�SCAND_MA�XyEI�c8�@FAIL_IMGy@�f���#�8�@IM�REGNUMyG
��KRSIZyC,����$,SONT�MOUW0{D�%��VU�#�c�� ��P�2FR:�\�O � �MC:\XS\LO�G�VB@4 !��O�_�Q�_o
�z? MCV�_�SoUD10fEX9k�
�f�wV�2ۜ�z�p(��=��͓o��j�o�o�o�o�o �o�o 2DVh�z��KPO64_r?S�0��n6�u�Q0LI Q�z�x�qV�� �|f@�w��w =	�xSZV�~w����wWAI���DSTAT ܄�;�@�_ď֏�$���EP12DWP�  ��P G�/����q�AP-��B_�JMPERR 1�ݜ�
  � 23�45678901 �������ʟ��ϟ� �$��H�;�l�_�q�x���LT@MLOW��8�P�@�P_TI_X�(�'�@MPHASOE  53���CSHIFTUB1=~k
 <���O b��A�g���w���ֿ ���������T�+� =ϊ�a�s��ϗϩ��� �����>��'�t�K��!��#ޛ:	VS�FT1�sV�@MN�� �5��4 �0���UA�  B8*���Ќ�0p����b�Ҫ��e@��ME*��{D�'���q��&%��!�M�$�~k���9@�$~�TDINGENDcXdHz�Ox@[O��aZ��S����.yE����G�� ��2����������RELE�y?w�^_�pVz�_ACTIV����H��0A �`�K��B#&��RD�p���
1YBOX ���-����2��D�190�.0.� 83���254���2�p�&��robot����   pxN g�pc�  �{�v�x���^$%ZABC�3�=,{�낆;-!/^/ E/W/i/{/�/�/�/�/ �/?�/6??/?l?!	ZAT����