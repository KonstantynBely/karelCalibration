��   ��A��*SYST�EM*��V7.7�077 2/6�/2013 A�   ��	��BIN_CFG_�T   X 	�$ENTRIES�  $Q0FUP?NG1F1O�2F2OPz ?C�NETG  �D�NSS* 8 }7 ABLED? �$IFACE_�NUM? $DBG_LEVEL��OM_NAME �!� ETH_�FLTR.� �$�   ��FTP_CTR�L. @� LOsG_8	CMO>�$DNLD_F�ILTE� � SUBDIRCAP"m� HO��NT.� 4� H�ZA?DDRTYP� A =H� NGTHph���z +LSP� D $ROB�OTIG cPEEyR�� MASKa�MRU~OMGDsEVlFRDM*��DIS���� TCPI�/ �3 $ARPSIyZoK_IPFp�W_MC-�F_�IN0FA~LAsSS�5HO_� �INFO��TEL� P�����R WORD � $ACCE�� LV�$TI�MEOUTuOR�T �ICEUmS�   �$O#  ����!���
��
� VIRTUAL�/�!'0 ��%
���F���F�� 22+5� '�� =��!�!j?�����; Ax?�5�=2~;�#"SHAR� 1>9  Pf?O(4OHO7OlO/O�O SO�OwO�O�O�O_�O 2_�OV__z_=_�_a_ s_�_�_�_�_o�_@o oovo9o�o]o�o�o �o�o�o<�o` #�G�k��� ��&��J��n�1� C���g�ȏ��쏯�� ӏ�F�	�j�-���Q� ��u����ן�ϟ0���7z _LIST �1�=x!1."k�09��j�1{��255.��r����05i�2p���� ������̯ަ3诂�@_�� �2�D�ަ4`����װ��������ަ5 ؿ��O����"�4�ަ6Pς���vψϚϬ�� �$��Q>�$ % =� .6+5U�o!�R��)��0H!�� ����rj3O_tpd��31 � >�!!KC� ����(�'6��!C� ;�����!GCON� ������Osmond���