��   3L�A��*SYST�EM*��V7.7�077 2/6�/2013 A�   ����UI_CONFI�G_T  d� )$NUM_M�ENUS  �9* NECTCR?ECOVER>C�COLOR_CR�R:EXTSTA�T��$DUMM�Y37CMEM_�LIMIR$D�BGLVL�PO�PUP_MASKx�zA  �]8�ODE�
9C�FOCA �40VCPS)C��g �
HAN� � T�IMEOU�PI�PESIZE ޝ MWIN�PA�NEMAP�  �� NU_FAV�B ?� 
$HL�P> _DIQ?<� mELEMV}#UR� h� So��$HMI�RO�'XW ADON�LY� �TOU�CH�PROO�MMO?$�A�LAR< �FIL�VEW�ENB�=!%bC -"U�SER6)FCTNV6)WI�� I* �_ED�h"R!_T�ITL� -"C_OORDF8" &�USTOM0 �t $} RT_OSPID��$C�$n*PAG� ?Z�DEVICE�)S�CREqEF����'N�@$FLA�G�@ �"USR�VI 1  < 	\� ;2�<1�PRI�m� A�� [0TRIP�"m��$$CLASS  ���|1���R��Rq0VIR�T_1z?�0'2 )��U�)�_p�R	 ��,��;���D�2�0�3�3�1��� , � � �?��
 �� �1<ONO`OrO�O�O�O 8O�O�O�O__'_ �OK_]_o_�_�_�_4_ �_�_�_�_o#o5o�_ Yoko}o�o�o�oBo�o �o�o1�oUg y����P�� 	��-�?��c�u��� ������L������)�;�M� TPTX��݈p����  sX���$�/softpar�t/genlin�k?help=/�md/tpmenu.dgO����� �؏C�U�g�y����� ,���ӯ���	���� ,�Q�c�u�������:��Ͽ����)���9���F�6�3S�($ÿ����nϧϒ������1�1���3a�(Y��?�����3�"� 1�5�2 �\�6 REC VED��i�{��wholemo�d.htm��si�ngl��dou�b��trip���brows ��+�|��0�B��f� x������f�P�߾��dev.s��lh$���<�1'�	tS� ��<��� �������������� 2[� �0s����� ��0pE W&{���]�V P���//,/>/ P/b/t/�/�/�/�/�/ �/�/??��.?(?V? h?z?�?�?�?�?�?�? �?
OO.O@OROdOvO �O�Oh�O�O�O__ /_A_S_e_w_r�_�_ |_�_�_�_���O=o 8oJo\o�o�o�o�o�o �o�o�o"4] Xj8?����� ����0�B�T�f� x���������ҏ��� �O1�C�U�g�y����� ����ӟ�_��	�؟� ?�Q�oo ������� ���ܯ� �)�$�6� H�q�l�~�������ƿ ���� �2�D�V� h�zόϞϰ������� ��
��.�@�R� ��� �߱����������� /�*�S�e�4�F��� d�v�\�������=� 8�J�\����������� ������"�B <j|����� ��0BTf x���|���/ /1/C/U/g/y/�/�/�/�/�/�/	?:��$UI_USERVIEW 1���R 
����J?\?�m {?�?�?�?�?�?�?O "O4OFOXO�?|O�O�O �O�Oo?�O�O�OgO0_ B_T_f_x__�_�_�_ �_�_�_�_o,o>oPo bo_oo�o�oo�o�o �o�o:L^p �%������o ����C�l�~��� ����W�؏���� � ÏD�V�h�z���7��� ����/���
��.�@� �d�v���������a� �����*�՟7�I� [�ͯ������̿޿�� ��&�8�J��nπ� �Ϥ϶�a�k�����Y� �4�F�X�j�|�ߠ� �������ߋ���0� B�T���a�s������ ���������,�>�P� b�t���)��������� ������#��^p ���I���  �6HZl~) 3��!��/ / 2/D/�h/z/�/�/�/ S/�/�/�/
??�(