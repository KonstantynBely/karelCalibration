��  ë�A��*SYST�EM*��V7.7�077 2/6�/2013 A�Q  �����ABSPOS_G�RP_T   � $PARA�M  �  �ALRM_�RECOV1   $ALMO�ENB��]ON�iI M_IF1� D $ENA�BLE k LA�ST_^  d�U�K}MAX�� $LDEBU�G@  
GPCOUPLED1� $[PP_P�ROCES0 � �1��URE�Q1 � $�SOFT; T_I�D�TOTAL_�EQ� $,N�O/PS_SPI�_INDE��$�DX�SCREE�N_NAME {�SIGNj���&PK_F�I� 	$TH{KY�PANE7�  	$DUM�MY12� �3��4�GRG_S�TR1 � �$TIT�$I��1&�$�$T�$5&6&7&8&9'0''��%!'�%5'1?'1*I'1S'1]'2h"GSBN_CFG1 � 8 $CNV_JNT_* ��DATA_CM�NT�!$FLA�GSL*CHEC�K��AT_CE�LLSETUP � P� HOM�E_IO� %�:3MACROF2R�EPRO8�DRUeNCD�i2SMp5�H UTOBACK}U0 � �	�DEVIC#TI\h�$DFD��ST�0B 3$INTERVAL��DISP_UNI�T��0_DO�6E{RR�9FR_Fa��INGRES��!Y0Q_�3t4C�_WA�4�12HGX�_D�#	 d �$CARD_E�XIST�$FSSB_TYPi�� CHKBD_S�E�5AGN G�� $SLOT_�NUMZ�APRE�V��G �1_E�DIT1
 � Uh1G=H0S?@�f%$EPY�$OPc �0L�ETE_OKzBU�S�P_CRyA�$�4�FAZ0LACIwY1KR�@k �1�COMMENy@$DGV]QP� h���AL*OU�B? , $�1V$1AB0~ OL�U=R"2CAM_;1� x�f$A�TTR��@0AN�N�@�IMG_H�EIGHyAcWI7DTH�VTCYU��0F_ASPE�CyA$M@EX�P;$� Mf�C�FcD X $�GR� � S!1U`BfPNFLIC`~d
�UIREs3��AO}MqWITCH}cJX`N.0S_d�SG0� � 
$WARNM'@f��@� sLI? �aNST� �CORN��1FL{TR�eTRAT@0�T�`  $ACC�1"p '|�'r�ORIkP�C�kRT�q0_SF� �!CHuGI1 [ �Tz`u3IPpTYPVD�@*2 �P�`�� 1zB*HD�SJ�* ��q2�v3�v4��v5�v6�v7�v8Z�v9� 
wpO�$ <� so�o�h�|s1�PO_MOR.� t 0E�v�NG�8`TBA� 5c���A������]@����ϋP��0Ѕ*��h�`�
P�@�2� �,p�J�,p_Rrrqo@+�J�/r/�J�JVq@�C�j��m�g��usp*o�CP_}0OF� �2  @� RO_����WaIT8C��N'OM_�0�1ەq3�dwpPcD !�;����hP���mCEXpG�0� F�<p%r
$TFx�J6F�D3ԐTO�3&@yU=0�� �YH�24�T1��E�� �e��f��f�>�0CPDBG;a� mk@$�PPU�3�f):��A��AX 1�dUN�$AI�3BUFuFvqᡎ�! |�`��`P�I��Pr�M�q�M~�䠁�Fr�SIMQS��G��Q�E������MC{�5 �$}1JB�`S��}1DEC�������ܴz� ě0CH�NS_EMP�r#$Gg�=Ǎ@_��q3�
p1_FP󔞡TCh�@`�b��q0�c}�y�G�� V�AԂ�!!���JR!0ԂSEGGFRA.pv 7aR��T_LIN�C��PCVF$������Y ���Q��)Bݲ��( '���f�e �S���Q��.0�p�B�8�A����SIZC����z�T��g������QRSINF3��p�� ��?�������؉����Lot��G�*�CRC�eFCCC�`+���T� h��mh�SbA��h�*��f��:�D�d�c��C��PTA����w@��L����EV���jF��_��F��N&�G�� �X������1i��! ��,��h#RGNP��0qF���R�}�D���2}�LEW�N��Hc6���C�K��vqRcDx �:�L��ou2���A6N:`Co�$LGp���B�1aP��s@�dWaA?@���~0R���d�ME%`��d�_RAs3dAZC���z�OkqFC�RH`X`�F�`��}��,�ADI;� 6b� ��@�`�p�`5cn�S�@�1�7a�AMP���PY$8CU�MwpU��iQU� $�P��C��CG1������DBOPXWO����pO$SK��2� wDBT TRL�1	 ��Q0Ti� �P��DJ�4LAY_C�AL�1R !'P1L	3&@�0ED�Q5'h�Q5'̡۱DB�2�1!�W�PR�'�qD1 0�1" �P�A$�q$�� �L�)#�/�#mpR�0$�/�$C�!%�/��$ENEqr�&��/�#d REp�"'�H �O)@7"$LF3#$�#xBП W;���FO[ _D0m�RO(@���u���j���3RIGGE�R�6PA%S���E�TURN�2RcMR-_��TU�`?�u0�EWM����GN�P��zBLA��E��/$$P#�CP� "��&@�Qk�C5D�mpD�A#�p4\1i�FGO_AWAY�2�MO��fQg ��DCS_(<�QIS ����c �C���A����B�t �Cn��A"�FW���D'NTV@��BVkQ��@���S˳W�sU�J&�xU�� ��SAFE��ZV_SV6bEXC�LUl�����ON�LA��SY��Q�tOyTBa��HI_V/>M�PPLY_�a��VRFY_#�q�B<d�_ )0��_+�Ip  �TSG3��b݀�0  AM���a*����0���Vi.b%fANNU�N� rLdIDp�U�2~S@�`mija�rj�f�pOGI:�"+��$FOb��׀OT@w1 ?$DUMMY���d�[!�d١�& �E,o ` 8�HEx�s��b�SB$�SU7FFI�@ (��@�a5�g6�b�wMSW�E- 8���KEYI����TM`Z1^ӌq�1�vIN��p���b. D��oHOST? !�r ���t[ �t٠�tYp�pcEM>���$���p�L��UL��/ p�|3��r�DT50~�!0 � $9��ESAMP�ԕF��������I�0��$SUBe�Q�� ��C�:��G�SAV ��r���G�C� ˇ�P�nfP$80E��YwN_B�1 0��DIad�@O���}�$]�R_I��� �ENC2_S�T � 2
ԇ J����L�q~S�`;����!3��M�I��1:�p�4  L�3�M��0��0K�4'a��AV�ER�q��}�M�DSP�v��PC�U����iì�VALU�ŗHE� ��M�I�P@���OPP7  ��THS ���6�SH�F�F􁳠dL��0�T��SC�Q�d�:�ETo�5zrF?ULL_DUY�da��0��O�w�h�OT��P���0NOAUkTO�!6�p$�H\���cl�
�C�P%�C�������L�� 7H *�L���n�b���$�0P�˴��ֲ��[!����a��Yq��dq��7*��8��9��0����U1��1��1��1ȺU1պ1�1�1���2
�2����2��2���2Ⱥ2պ2�2��2��3
�3��3T����3��3Ⱥ3պU3�3�3��4
��Z���SE�"8 < ��~��`�;I�����/��QFE�0�0� �9 ,��Q? z@^ ?�А��ER@#��Q�A��z� :�`$TP�?$VARI�<�n��UP2�P; �pq�TD��S|�1`3�p���`!r�BAC�G< T�pr��)�p�bP�P o�IFI)� P ���U���P��P���0��� =t �;'�Ԡ��P'�ST (&�� HR&�r0E��*��	%�C��	��� _Cr�N�r��B��p�h�FORCEUP%b^n�FLUS�`H�N �E�h�RD_C�MK@E(����IN�_��&vPg�REMM�F~Q��M �� �3
K	N0�EcFF��N@IN�A��OVMl	OVA�l	TROV���DyT��mDTMX� ��m{@�
��? �*X[ ��CL��_:p�']@$�-	_
�;_QT��X
��@AQ	D� ��}��}!�V1� RQ��LI�MIT_�a椀�M���CLmd}�RIqV	�a��EAR��IO*PCC�����B�Bg�CM@��R{ �GCLF��G!DYM(/�aR#5TWDG��| s%�Z�FSS& �s> �P�a�!r1��wP_(�!�(�!1��E�3�!�3�+5�&�GRA����?w��kPW晅ONT��EBU�G)S&2*[�{@a�_/E @�P�Q3�_�TERMB5AK5���ORIG0B<K5���SM_�Pr�rG0CK5g@�TA�9�Dd6[�UPB�Eg� -zAa�@.P|Y3.@A$SEG�:vf ELEUUSE�@NFI,��2�1xޠp4�4B$UF6P�$�FQ4@�wAG0TQ�&�HSwNST PATm�<piBPTHJ�AߠE�p��2�P؀	E)��؁��1R�@�InaS�HFT_��1oA�H_�SHOR ܣ�6 ��0$�7�@Dq�'�O#VR#�na�@I�@��U�b �QAYLO=�z��I'"�oAj�!�j�ERV��:Qh� �J��OG @�B0����U�>���R!P"�AScYM.�"��1WJG�уES�A�YvR�U�T @���E)�ᥳEaP!�WP!�WOR @�MB��GRSMT�F�GR��3la�PA.@��[��q�uG� � ����T�OC�1�`P�@ �$OP��ဝpՓá� ��O��RE�`RC�AO�pтpBe�`RmE u�h�A���e$PWR�IM�ekRR_�c���q.B H2H���p�_ADDR��H_LENGqByqnq�q��R��S�I H��S���q0Ӧu>Ӵu���u��SE�'�LryS��J $�<�`��_OFF��r�PRM� ��aTTP_�H��K (^pOBJ�?"ip��$��LE�`C!�ȠL � ��׬�AB_~T�S�s�S{`��*�LV�N�KR��eHIT���BG��LO�q t�fN�͂���`���`3SS{ ��HW��A��M�p`INC�PU�"VISIO �����+��t,��t,�~�� �IOLN���N̠�C��$�SLQb��PUTM_�$�`{�P x�V���F_AS�"O��$L��I���D�A��U�0�@Af��`q�<PHY���Ó�;ថUO��#P `������ڔ� �2�pP���`(�L��XY�B���UJ�Q�vz�NEWJOG-GN��DISx�[�K-�Lf�#R 
�WAV��ǢCTR�CǢFL�AG�"[�LG�dS� ���Y�3LG_SIZo�����X����FD)�I� 4�E�*��D0���c $���𖶦���K���xD0��� SCH_���߅p�2��N��F�T
���E�"~�����"��U
�
�{`L�	�7DAU/�EA�-�؞dE�;�GH�b<*����BOO��U�h Aɒ��ITp��y�[0ŖREC���SCR��ʑDI2ēS.@��RGO����˒����d�´���S�U���W�Ĳ�Ľ�J{GM$�MNCH,󾲑FNKEY%�KnM�PRGK�UFY��PY�FWDY�HL.��STPY�VY�@XY؀�Y�RS��H1`uۺ�CT���R��� �$�U	�m���
R��ݠғ`�G=��@PO�d�ڻŦ�M�FO{CUd�RGEX���TUIK�I{��� ��	������I�M��@A�S�`���@������ANA���2�V7AILl�CL!�U?DCS_HI+4`�D�s_�Oe�
!h�S���|�S����IGN 4��F�J��T�b�8�BUj � V !PT�$*��rvP�Ϥ�!��AVrW �!Pi�'���0�1
?2?3?t���`�>� X � i�=a0�5���Ņ�ID� tb	P5R�bOh ��\A�+ST	�RF�Y� �@~�  W$E�C�y�������!Y L�؟0� �@���`qFtǀ�Fw�Ҭ�_ Z ��p����b���>0C���[ �p CLD�P	��UTRQLI�{��T����FLG �� 1�O�D������LD���ORG������hW>(�spiT�r� 4\ �#0P��վ�Sy`T��0#0' �$�!�#RCLMC�$B/T/�)�Q��!=1I�p_d] �d�RQ73$DgSTB�p�   6l��-8AX�R /8>I<EXCES�b�R2Mp�1^�p2��T�12��0_�p"6_A:&��;G?Y8�0K�d` \�G�ROU��t$MB� �LI9�CREQGUIRDB�aLO#KODEBUr� 1LYM��agb��`@�C6�"0ND��`�c`b���̨�CDC���IN'��C��Z`���H��N��a#�� � 1�APST�� �c\rLOC�R!ITp��P�Ap��1 1ODAQ��d� X��ON�cF �R�fV�	X��b�U����uFX0IG}G�� e �y @X�a��X�XR�Q%��Y	��X	��V<�0ғDATA$`�E�a��a�N��f t $MDEaI:�)Sf��^d�![g�H5P�@]ez��a_cANSW�a^d�a��^e�D�)ARz�� Xpg[ �0CU4�V�`��=URR2{�h �D2�`A��A�! ?d$CALI&0���GS�w2K�RINtb�t<�NTEg�(i�bCu��=RBqg�_N�qjPukr���$tht�2kuyDIV�&�DHi0jp+�l c$Vp�C�$M�$Z�<!T �����b�emH ��$BELT˪ZA/CCEL���;�"�IRCO�݁m��yT���$PSi0
�L�0ڰW��Cp�8��T�9�PATH���.���3]��Pl1�_<�r��Ł�"S C�r��_MG��$�DD�9���$FW�`7`���.����DE�PPABN�e�ROTSPEEՂ@L� JN�@���(0��0$USE�_p�P&�ܦSYh>��p�! �QYN09A����OFFua��7MOU߁NGJ�܀sOL~�ٔINC�d�2Q��-2��� -2ENCSpa2U��,+4R�IN�I]�B����"n�VE��s^��23_UPօp�LOWL��[�` '���D>�2@Ep]�'��2C[pW�MOS����4MO��0�'P�ERCH  ��OV����蓼����� �$�8S+�� 2@����B��V�0^�O�L�0P��7O�U�UP"��������TRK��AYLOA�J��1���]�͵³3P� �RT1I�1	�� MO�_��-2�28 �`4�w�ٳ��?�pDUM2���S_BCKLSH_C]�P�ϐΦ� ���bn�"�y�Ñ��!CLAL V��!���� ��CHK �SՐRTY����C�
�*!6a_�ä_UM�����C���SCL��W�LMT_J1_L< 0-օa:�E4�U�G�D�J�P�J�SPCd�ȑZ���3�PC �3�H_A@�2��C� cXT���CN_rN���.�S��%�V���:� ���]�9���C' �SH�r�*�*!9��9� p��^���9���P�A���_P��_ �"�Ŷ�!ճ����cJG����~�OG�׾,�TORQU��ON��޹*�B٢-�*�&L�_Wž�_�sj�P�sj��sj�Ir�I��%I�sFKP]�J�!��,c!�VC�0'42���1��{0��82��J�RK��+� DBOL_SM���"M�@�_DL�q�"GRV�q�j�sj�sKH_p��I���
COS��LN- ���� �p�	�p�	�����bFZ� ٦KMY��D�TH�eTH�ET0��NK23��s��s� CB�CB�sC&1n2�����s��SB�s��'GTS�1W�C.�2Q������$�'3$DU���8A!r��2P&�1Qb8V$NE�4�PI� ���"$%�v$�p�A��%p�'���LPH�5�"h��"S��3�3�3�"+3:2�pV��(V�(�p�,V�*V�;V;V";V0;V
>;VL9H�(�&�2�-�n�H;H;H";H�0;H>;HL9O�,OR�(O}I�.O�*O;UO;O";O0;O>;O2F�"�Y�T��'SPBALANgCE_T@SLE�H_�SPHq�hR��hR3PFULC�lX�R{W�R3Uz1i�
�UTO_����Tg1T2�Y�2N�� �`��Tq���Ps d���T�O�p!�L�INSEG���R�EVf��Q�DIF̨�zy1j_g�r1k���OBUa��t$yM�I`���SLCHW3AR>��AB��u?$MECH�TXˑ�a��AX˱Py�p�f�'�r�Pl 
�b�I��:�ROB�C�RW�-u��:*��MSK_KP�tn WP �P_��R��r_tn���18�c�a�`_p`�y�_p�aIN:a��MTCOM_�C���po  �݀g`4�$NOR�ES��r��`�rp� 8U�GRJ��eS�D� ABג$XYZ_DA�!F�r�DEBU:a�q���p�q _P$��COD��� 1����`���$BUFIN�DXa�  !�M{ORRsr $�q�U&���u��ӑy�]�_��bGi�s �� $SIMUL���8��>���F�OB�JEjP��ADJUySψAY_I���8�D���s�Ԑ_F-Iב=s�TZ�� c����`b�"�(�b`tp0G�D��FRIWÚd�Tg�RO%�A�E�b񊰃^�OPWO�> Vpt0>�SY�SBU0[�$SO!P��I�����U��b`�PRUN�rڕPA�rpDٖ�b��1�_O�UTΑ�a�t$^�IMAG��\p�v PDaIM��1�I�N[ �0�RGOVCRDY�˒���P�/�a�� L_�PB�}�L���RB�� �љMkᜪEDb��` J�N�@M��~�w���]�SLjPVpu x $OVSLfwSDI��DEX��@�q�����o��Vb��N�A��'��,��'�D�M~Ҥ_�SETK�Vpv @0U�^��ep�RI��j��
q�_�}������^�dà*� w �H\q�`��ATUS><�$TRCx T��X�ѳBTMڷıI
��P�4}Ѱ���Vpx D\pE���β�0Ehbϱ�����ϱEXEհ����)�=���f�ym�]p԰UP��L�$�`6�XN�N���������� ��PG�uzWU�Bñ�e��ñ��JM/PWAI[�P��œLO7��pFA`���$RCVFAIL#_Cwq�p��R9��p��c��(�}�"�-�AR�_PL��DBTB8��,��pBWD ��p3UM*�"�IG�7��Qc�TNLW�"�}�Ry�iӻ�E�����|����DEFSP` { L\p�`��q_��Ճ��UNI�����Ѐ�RD��Rb _ULA`Pͱ��P�pUq|-�#��q�O��tXPc�N�PKET��
��Pq�Uq} �h�ARSIZE�5p��=��u�S̀O�R��FORMAT��Pg�COנq�<bEeM�d����UX���,�Z�PLIb�Uq~�  $�pP_SWI�`V�/ G�b�?AL_ o��ХA�rB���C�rDn��$EL����C_lі� � �� ���r��J3x0 �r��TIA4Z�u5Z�6�rMOM��@f��s���pB���ADf��s����PU�NR����s�������Rt�� A$PI�&E�kqE� p-~-�-�W@C�0$��&�9q��gE��eSPEEDL@G�����Ծ�� ��)�9����)��	)���SAMWPx�08�1��MOVD�H$�_S`Y%nk%_��1�t�2�t����c�vd��8�H�PxIN� ��������(x�+(+GAMM<V|u!�$GETE��U�ٓD5��r
�PL�IBRv���I�$HIu�_L�ݰpB�&�E�(A�.� �&LW�-�&�,�)	6�&1���f�`j��� $PDCK���ٓ_���r�E��ီb7��a4��a9�� _$I��R�`�D�c�b~�Ե`LE��qkq���81��0�6pHp��`Vp�P/a?UR_SCR��A��r��S_SAVEc_D��8Ex�NO5�C��y�6�8@{$E�. {I��G	{I�@�J�KP �q��H� ���x" Mao���s���� d��6W2U�Cqy�ѡ:��M� �k�F� �aE��3�W<�@[�BjQWg@5r�U�R�R���Sc2jQM"��[C�L�W��M)ATr� ?� $PY����g$W`�fNG� O�`�b�b�b #�HЈ��a� ���c��%X�O���Z�e��ހRt� p䠰p�3+zO�O�O�O�O�a:5�_�r� |�E� 8@��>vs�>v��8@_��kwVvy�Eހu% Q��"rB�\�P�"tP���PM&�Q}U5 � 8*��QCOU�1 �QT�H#pHOL<�QH�YS��ESe�qU�E�p.BZ�O�� � q�P���%��UN\ְ�Q ��OE��p� P2�3��AÔ�ROG�����Q2(�O}�2�������INFO�q� �#�e����RȾ�OI� (�0SLEQ�с�рi�C�{�ID��L��`� OK0�r��!E� NU�!��AUTTA�COPYqu�?��`@EML�NI�M�X�C���� Y�RGADJʵq�i�X�Q��$Pഖ�`��W��P��`�0�������EX8�KYC0b�Obpr�q���$�_NA9!�������`��?� � Q����POR�A�B�S�RV0�)a�Y�DI��T_��{������P�������5��6��%7��8y��S8BL�=�m�MC_F�p��PL9A8An�ȰR ��9��Ѽ��$iB�����d� ,�0FL�-`L�C@YN�[�Mz��C?��PWRc���L��!�DELA���8Y5�AD�a��qQSKIP�� �Q�4�OR`NT2�Q ��P_4�� ַ@lbYp�� ��������Ƞ��ՠ���������9�1��J2R� L�� 46*�EXs TQ%�� ��(Q����p�����p��̀RDCf� �`��X9�R�p������r��A$RGEA�R_� IOT�2F�LG��vi��M%PC���B�UM_����J�2TH2N'�� �1�����G8 TN00 �����Ml��`I�8eQREF:r1�q� l�h���ENAB{�(cTPE�0�1���i�m� ��^QB#��:��"������2�ҙ������P����&�3�Қ7�@I�[�m���&�4��������������&�5�Ҝ1�C�U�g�y���&�6�ҝ������P����&�7�Ҟ+@=Oas�&�8��������&�SMSK�q�|��a��E?A��MOT-EF����a@���(Q�IOQ5�Itc(P��POW�0L�� �pZ�����#p%�L��U�"$DSB_SIGN�1�)Q%���Cl�(P�P�_RS232��b��iDEVICEU�S�,R'RPARI�T��D!OPBIT�`QY�OWCON�TR;�(Q��O'RC�U� MDSUXTA�SKT3N�p[0�$T�ATU`P�S��0L����p_,PC�9�$FREEF�ROMSp��%�GsET�0�UPD(��A�2�#P� J���� !)$US�A^���6���ERcIO�P@bpRY�5:"_>@ �P}1�!�6'WRKI[D���6���aFRIEND<mQ�P$UFw����0TOOLFMY��t$LENGT�H_VTl�FIR��`-C�RSEN ;IU�FINR]��R�GI�1ӐAITI���4GXӱCI�FG2�7G1��Ѐ3�B�GcPR� A�O_~ +0!�1REЀ�E3�e�TC���Q�AVG �G8��"J���u1~! ��J�8�%���%m��5�0G4��X _0)�L|�T�3H6��8���%r4E3%GU�W�P�W�R�TD����T��а��Q��Tm�$V 2!����1���91�8�0U2�;2/k3�;3�: iva�9=i�aa�^SL�jR$V��SBV�E�V'�V�BK���� �&c�p��F�"{�@��2q�PS�E���$.rRC��o$AŠFwPR��Gv]U�c�S'�� 7�?8I�� 0�@qV`��p�d`A���E0�@��=�
B5�S!� ��aRHg����R�6�N SAX�!$�A�0L(A����rTHIC�1pY���h�t1TFEI�|�q�uIF_CH�3��qI�G�a�pG1@bxf���m���S@��7_JF��PR�ֱ��S��Ԁ�d ӎ$SР�Z�GRsOU�̃TOT�t�̃DSP�JOG����#��_P��"O������j��&KEPF(�IR����@M�R&@�AP�Qn�E^�`�!�[�SYS6��"[�;PGu�BRK�B �.��pIq�p��M���΂�`AD�!̃9�OBSOC׆�NӕDUMMY14�p�@SV�PDE_O�P�#SFSPD_WOVR=���C�L��OR�CNm0b�F.����OV��CSFR��pU���Fn���!#��C��A�"LC1H����РOV�s0���W�@M��ĥ:�R�O�#ߑ�_�p��s @@�u@VER�pns0OFSu@CV? �2WD6���2�ߑj2,Y���TR�!����E_FDOY�MB�_CM�D�B�BAL�b>�f��attV"Q �240/p��N�Gg�z�AMx�Z�0���¿�_M~��"7����8�$CA�7�D�����HBK81��I�O�5���QPPA�=�"�M�5�͵�~��DVC_DBxC�~� �3"�Т�!��1��糖�3����pЈ��*��U�3��CAB��2VӆPѣIP���c�O��UX�S�UBCPU�r	�S �P P���90^SQ׹c���."��$HW_AC�Т��S��cA�A~�pl$UNIT��}l��ATTRI"����	�CYCL��N�ECA��J�FLT?R_2_FI_�G(��9&�1LP�?�>�o_SCT�CF_��cF_��6��FS8!����CHA�1�w�8���"v�RSD�4"�����q�_T��PcRO��>�� EMy�_ܠ��8d��a 1d��a��DIb0!�?RAILAC��9RM��LOÐ C��Q�*q��3q���PRJ��SQ�pU�Cr�zs 	�FUNC��@rRIN'PѸ0���u��!RA��B �����F�Ğ�WAR�~���BLQ����A0��������DA����	����LD)0��Q�1�q��*q1TI�2rQǁ�p$xPR�IA1�"AFB�P�!|ߠ�<`�R����MOI��A�DFa_&@��51��LM��{FA�@HRDY�4ORG6 H���A�0| �MULSE&@x"�Q��a �G��	�����$dm$�1$1 ��|�0���� xm��EG�̃�`ARހ��09�2o���z�AXE�ROB��W�A��_�œS�Y������S�W�RI�@s1��SCTR�� ��(�E�ч 	%1��AB�( �/&�a�ӰOT�0^�	$ߠARAY�sf"���S@	��FI��*�$LI�NK���!�a_�%#�%{q�"X�YZ82�*�q�#OFIF���"�"�(j 	B�j�4С��n�3FI��%7�q���j���_J���%��#N�QOP_>$H+5�3F�PTB\1�2C�Цi�DU�&62�TURN��2r�5t!}��p��|7FL�`��Ӑm�0�%+*7�	� W1�. K�M��&82�Q�2rQ�#�ORQ��G��-(�+p���z�� 3q�E"��TF�GOV�@-A��M*��y�4�E:�E@�FW �J��G���D��o�*� � ��A7�P��y��E��A�GZU:ZU�CG�E)R���	6�E���B�TAFQ��)4����0r'�AXУa2 .q�c�W�c�W�c�W �p�Z�0�Z�0�Z%@�Z K@�Z��Z
!�V� �Y � 
i� i� *i� :i � Ji� Zi� ji� zi��a�iDEBU{�$v�u��;q��"F7O�n�AB��6��C9V�z� 
fr�� ��ukњw�!�w�!�w �1�w�1�w%A�wKA�w���\0��"3LAB"2|EwЄ�҂�3� .*�SE�RVEN� �� $q�_NAǁ!_�PO����` xf�EP�_MRA��_� d  T�����ERR����~ T)Yi��RI�V"0�SN��TOQ�T)PL��T�Ѕ ����J_ � p�PTl X���_V1�b�Q���#�2�2+������/@��p��5�$W���V���VN�[�$�@�� �S���Q��	EHELL_C�FGN� 5�%�B_BAS��SqRvp0�K� �QS��Jϐ1a�%ΑU2�3�4�5�6�7�8�RaO���� � NL:Ɵ3ABn��АACKwv��)�o�u0�iႩ_PU2�CO,q��OU��P��ӕ`�����TP��_KAR�0��R�Em�� P����Q�UE٩��@���C�STOPI_AL zs��� �TĠ�� GSEM[�w�k�Mw�6y�TY��SO`��DI���Є�=�װ�_TMK�MANR�Qζ� E��$�KEYSWITCaH��Ѱ��HE��OBEAT���Ep�LE����&�U��F�d�����SO_HOuM� O��REF�@�PRi��R� ��Cr@�O0�p ECO��|�� _IOCM�4�M�k�K���'�O�# D�!ۧH�U��;��M7��@�3FOR9Cߣ�� q�����OMq � @�Etxk�U#Po1(B�O�o3B�4x�NPX_AS���; 0ݐADD��(��$SIZߡ$�VAR�TIPRr�q�G�A(ҷ��@
�˨r�t�n�SV��XC����FRIF��R��S%�7�x���N�FѲEАO� x6�PSIڂTEC*�.%CSGL=�T�"�0�&�V�D��>�ST�MT
�o�P\�ByW�@?�SHOWw���P�SV� K�w� ���A00�0 �Q��K���O���_���Ti���5��6��7��8��9��A����@6���������F�� 
 ����U ����� �����0�� �J@��:�1�G�1T�1a�1n�1�{�1��2��2��2���2��2��2�2��2 �2-�2:�2�G�2T�2a�2n�2�{�2��3��3��3���3��3��3�3��3 �3-�3:�3�G�3T�3a�3n�3�{�3��454��4���4��4��4�4��4 �4-�4:�4�G�4T�4a�4n�4�{�4��555��5���5��5��5�5��5 �5-�5:�5�G�5T�5a�5n�5�{�5��656��6���6��6��6�6��6 �6-�6:�6�G�6T�6a�6n�6�{�6��757��7���7��7��7�7��7 �7-�7:�7�G�7T�7a�7n�7�{�7��K�VP$�U�PD��  ��P���x�YSLO>��� � ��հ0�����QTAS�sTƠ��ALU}U�����CU��WFdQID�_Lѳ�UHI�ZI~�$FILE_Σ��T�$u�_VSA΁�� h��+`E_BLCK(�8bg�AhD_CPUQi��Qi����Sod_R1�ɢRw ��
PW,�d� �aLA�Sp���c�a�dRUN5� �a�d�a�d��5��a�d��a�d �T�pAC�C���X -$&qLEN~�3t���&p����Iѱ
�LO�W_AXI(�F1&q�T2mwM��ɢ�����I����Q�yT#OR.�&p�{DW��s�LACE���&p8�����_MAuйv8�u�w�qTCV�|��wTڱ�;�1�<ѷt���_��s��J����MD��ӠJ����u��
�u2q2�������l�s�pJKцVK~�hか��3ՃJ0����JJ�JJ��A�AL�����42�5Xr;�N1B�N�(�	��tL�p_k��x��"p��� `5`�GROU�PY�ӲB>$�NFLIC�ө�REQUIREv�EBUV�"q���кp2���#pɖ!qxг��� \��APP�RՐC���p
!�E�N�CLOz�,�SC_M ���A��u
!q޸�� 䣠MCp�r;�Xr|�_MG���C��,`��N��p��wBRK��NOL��t����Rϰ_LI��Hէ����JޠѤP� �p��p���p;��pD�"�p6�K��8��n�|"q���� Ғ�Mr:ql�Gqz�PATHv�������Rx��������pCNR�CaA��է���IN%r�UC�pwQ�Cd�U�M�Yop�����QE�:p�Gp�����PA�YLOAͧJ2L�HPR_ANqQ�L��`[�W�K�g���R_?F2LSHRё�LO\�䱕����ACRL_������޷C�XrH�P"�$yH���FLEX�� qJ%u� :2Dv�p4�K�GYq0�pPbt|F1Kљ� �׃�������E����/�A�S� e�w�����y���ф��@�蘏����J�ÊT���X����υ ��څ ��[����
�� �)�@�;�D�V�h�z��>��� � �������QIPAT��ё���EL4� �ؘJڿ��ߐJE��CTYRޱ��TN��F��ɗHAND_VB�p�ѹP`�� $�&�F2��K��ШRS�W9 qj��� '$$M��}�R��E@��Uw�H��sA�P H����Q���A���P
��A��Aɫ���j`���D��DɫP��G�`1)ST��9!��9!N̨DY�`���| �Y�鰋�KыǦ�J� ч�s�U�ХP���&�/�8�A�J�S�Y�J��� ; �t�.Rx66N�/QASYM����Ґ����Խ��ٿ_SH�����筀�4��+�=�O�J�V��h�'CI����_�VI�dHN�u@V_UNI�ÉD���J҅�B�%�B�̦D�� �D�F�̓��������$*Uc���Q=��H�`��XQE�N� v�DIɠS�O�wToY�YP��� ��I�1A�Q�äQ �`Bc�S`�  p�a.a�� � MEB����R'RDaTkPPT�0) ���Qz�~�A��0�Xa	iT@�� $DUM�MY1��$PSm_��RF��  ���Pf�aLA��YP��jb�S$GLB_T>mU�e�PpQ p8���Q� X	�ɗ�`�ST��ߐSB}R��M21_V��8$SV_ER��1OÐ�c�cCL�`�bEA5�O�RTPT O�P � D �`3OB���LO˰&u�q9c�`r�0�SYSqADR�TP�P�TCHb � �,&����W_NA����tz���Y�S�R���l  =��M�u`�ys�u ~�s��s����� ������0�)�T� "�5�~���B����s�?��?�?DY�XSCR�E)�p�ȐST[�s}�P!��t�QQr _� Aq� T	��`ob��a`��l��Ҥ��g�c�O�� IS�c��TuvY�UE�T� �ñ�jp^`Sq�RSM�_iqmUUNEXCcEPlV֑XPS_�a ����޳����޳R��COU�ҒS� [1�d�UE�tҘR|�b9�PROGM� {FL�$CU�`cPO?Q�д�I_�P}H�� � 8�.��_HEP����~�PRY ?��`�Ab_�?dGb��OUS>�� � @�`v�$BUTT�R|V`��COLUM�<�U3�SERVx��OPANE� q��P�@GEU�<�F����q)$HELP�B�l2ETER��) _��m�Am���l����l�0l�0l�0Q�I)Nf��S@N0�� �ǧ1����ޠ ��)�LNkr� Ʉ�`T�_B���$9H�b TEX�*�x�ja>�RELV�СDIP>�P�"�M�M3�?,i�0ðN�ja�e���USRVI;EWq� <�`�PuU�PNFI� ���FOCUP��PRIa0m@`(Q���TRIPzqm�sUNP�T� f0<��mUWARNlU��_SRTOL�u����3�O�3ORNN3�RAU�6�TK��vw�VI͑�U�� $V�PATyH��V�CACH��LOG�נ�LIM��B���xv��HO;ST�r!�R��=R<�OBOT�s��+IM�� gdSX`} �2����a���a��VC�PU_AVAIL�eb��EX��!W1N ��=�>f1?e1?e1� n�S���P$BACKLAS��pu�n���p�  fP�C�3�@$TO�OL�t$n�_JM�Pd� ݽ��U�$SS�C6X`�V�SHIF ��S�AP`V��tĐG�R+�^P�OSUR�W�P�RADI��P�_ cb���|a�Qzr|��LU�A$OUT?PUT_BMc�J�IM���2��=@zr��wTIL��SCOL���C����ҭ�Һ� ���������o�od!5�?��Ȧ2Ƣ)�VVp�U���vyDJ�U2Ѭ�� �WAIETU����n���%��{NE>u�YBO�� �� $�UPvtfaSB�	TPE/�NEC���  �ؐ�`0�R6�( �Q��� ش�SBL�TM[���q��9p����.p�OP��MAS�f�_DO�rdATZpD�J����Zp��DELAYng�JOذ��q�3�����v0��vx��,d9pY_ ���	�7"\��цrP�? �QZABC�u� ��c"��z��
s �$$C��>�����!X`xs � � VIRT����/� ABSf�u�1� �%� < �! �/�/??0?B?T?f? x?�?�?�?�?�?�?�? OO,O>OPObOtO�O �O�O�O�O�O�O__ (_:_L_^_p_�_�_�_ �_�_�_�_ oo$o6o HoZolo~o�o�o�o�o��o�o�o{� ��AXgLMT�s��#7  �tIN&8q�tPREO��+v�upXuLARMRE?COV �)Xr�zujF �%/�!d� �����7�I�[�<m�~�, 
�/���vNG5� �+	? A   ڏ싾� PPLIC5�?��%upՁ�Handling�Tool -� �
V7.70P/�36뀬�
]�_3SW2�D�F0j�W� 43Y�J�9�K��7DA7?�����
&�X�e	-�N�one��J������ �T7�	���_�Viu�6s��UTOz"�,t�Ty.�HGAPONЬ %��!.�U��D ;1�y� t�x������y.�K�Q 1M�{  Hp������	���uq��"��" ��!��Hեw��?HTTHKY��" ٯ����u������ ��Ͽ�����)�;� M�_�qσϕ��Ϲ��� ������%�7�I�[� m�ߑ��ߵ������� ���!�3�E�W�i�{� �������������� �/�A�S�e�w����� ����������+ =Oas���� ���'9K ]o������ ��/#/5/G/Y/k/ }/�/�/�/�/�/�/�/ ??1?C?U?g?y?�? �?�?�?�?�?�?	OO -O?OQOcOuO�O�O�O`�O�O�O���TOĀ���DO_CLE�AND���{SNM  ɋ���_�_�_��_o��_DSPDgRYR�_��HI!��]@�_}o�o�o�o�o �o�o�o1CU��MAX �bTQNQS�sqXbTB�o�B���PLUGGb�cWo���PRC4`B�P"]klo^�rO�r=o^��SEGF;�K� +�6��_�_}�������8ŏ�0�LAPZom� /��+�=�O�a�s����������͟ߟ�6�T�OTAL�v�y6�U�SENUZ�g� �HXL�NR��RG_S�TRING 1~3�
�M,��S�
��_ITwEM1��  n� ����Я�����*� <�N�`�r����������̿޿��I/�O SIGNAL���Tryou�t Mode���InpB�Simu�lated��O�utT�OVE�RRW` = 10�0��In cy�clHŕ�Pro?g Abor^Õ��>�Status���	Heartb�eat��MH �Faul����Aler�����'�9��K�]�o߁ߓߥ� ^S��^Q������� �,�>�P�b�t��� �����������(�:���WOR9���r� ��L������������� *<N`r��������PO�������9K ]o������ ��/#/5/G/Y/k/8}/�/DEV�  -�/�/�/??)?;? M?_?q?�?�?�?�?�?��?�?OO%O7OPALT��^A��8O�O �O�O�O�O�O�O__ (_:_L_^_p_�_�_�_8�_�_LOGRIxp�� avO�_*o<oNo`oro �o�o�o�o�o�o�o &8J\n�_*�R�ݦqo���� ��(�:�L�^�p��� ������ʏ܏� ���PREGbNK�� $�r���������̟ޟ ���&�8�J�\�n������������$A�RG_r�D ?	��������  	]$�	[�]����.��SBN_�CONFIG ���L�K�F�C�II_SAVE � �k�b��T�CELLSETU�P ��%  ?OME_IO��%MOV_H��¿ȿREP�|��UTOBACK���V�FRwA:\8� �,8���'`��8�cϮ,�INIa@8��^�,�MESSA�Gz��������OD�E_D��}�C���Ox� ��,�PAUS�!��� ((O��J�\�F�|�jߠ� ���߲����������B�0�f�t�%�*TSK  5ݒϕ�/��UPDT����d�����XSCRDCoFG 1���' �������&� 8�J�\�n���\�n�� ��������"��F ��j|����/�e�2�GROUN�����UP_NA�ܰ��	2��_�ED��1
��
 ��%-BCKEDT-��}��pg�Hg3�p8�e/�/�8���gA2���E/��/���/~/��ED3 n/&/�/J/\.�/"?�/�/ED4?�/?�/�\.[?�?5?G?ED5 �?n?#O�?\.�?jO�?�?ED6ZOO�O6O�\.�O_}O�OED7 �O�Ok_�O\.G_�_!_3_ED8�_�o��]-�_Vo�_�_ED!9Fo�_�o"o]-�o�oio{oCRoY_V h�]1�{� L?NO_DEL�GE_UNUSE�	LAL_OU�T V��W?D_ABOR���~��5�ITR_RT�N�ǀH�NONS�)Ю�����CAM�_PARAM 1�����
 8
�SONY XC-�56 23456�7890Y �~f�@���?�W�( А��8�h��х�ڎ��HR5pǃ��	��R570�B�Affފ��� ���ڟ�ǟ�"��� F�X�3�|���i���į�!�CE_RIA_UI������F��3;�Я ����GP 1���s�����V�IC󠸾����CO��C ��(��ǀC8ʺ�@��H��CCX�����Ch��p��x����� C�����Ⱥ��+�=�G���ށ��HE/pONF�IG=�f�G_PR/I 1�B�$ r����������(��~�CHKPAUS�� 1���� , wuj�|ߎߠ߲����� ������0�B�T�f�x����D�O����T��_MOR�GRP 2?� y�\�� 	 � ,��P�>�t�b���5�"����e�.�?a�a������K���d�P��V��a�A-`�/A�

 s�������b&��i��ܦPDB������)
mc:c?pmidbg���:�  g������p�U �  ����pM�3� ��d�/  ��{C��e�/��/��b{g�+/� O��}f/s/i�u/�
?DEF �(K��)�b buf.�txt�/�/��_�MC�����d(,53����ʇ��Cz  B�p�B��5�Bma�B�!)BR�Bs�UB��
�q�Dv��C��C���D"L�D;�ZD��:�=F��F�|ḚZFn�ߊF�2?E����_�:����S4���(D~���/��ʄ3@�à1/  TB�D=�V@a  EI�5�� F*� F��G$ˀF[�� GR��<Gl���G��G���&H��G֓ϦH���8b�� � >�33 9�ށ�  n^���@߂5Y�Ed��A���=L��<#�
 ��_�*~2RSMOFS���.^�9T1��D�E ��l 
� Q�;�P  x0_*_>TEST�")__��R���#o�^6C@A�KY���Qo2I��B���� �C�qeT�pFPROG %�(S�o�gI�qRu�����dKEY_TBL�  6��y� �	�
�� !�"#$%&'()�*+,-./01���:;<=>?@�ABC� GHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~�����������������������������������������������������������������������������q��͓���������������������������������耇���������������������9�Eъ`LCK�l��<�`�`STAT�c_AUTO_DN ��O�INDTO_ENB;���R�Q�Y�K�T2����STqO�~��TRL�`�LETE�ފ_�SCREEN �jkcsc� 	�UπMME�NU 1i  <�l�ol� K�u���FS����柽� ϟ���R�)�;�a� ��q���Я�����ݯ ��N�%�7���[�m� ������ɿ�ٿ�8� �!�n�E�W�}϶ύ� ��������"����1� j�A�Sߠ�w߉��߭� ��������T�+�=� ��a�s������� ����>��'�M���]� o��������������:#p)+�_M�ANUAvՏ�$�DBCOu�RIG��$�DBNUMLIIz��,1e
��PXWORK 1k�_-<_N�`r�TB_� � m��Y0�_�AWAY��QG�@b=�P�_AL� =���YҀ��`��_�  1!�[/ , 

:&dP2/o/�&�Mt�IZP��@P�#ONTImM��d��&��
�e#MOTN�END�o$REC�ORD 1'k8U2)?��O�?1-? &k�k?}?�?�?88�? �???�?c?O*O<O�? �?rO�?�OO�O�O�O �O�O_�O8_�O\_n_ �_�__�_%_�_I_�_ o"o4o�_Xo�_|o�_ �o�o�o�oEo�oio �oBTfx�o� �/�����>� )�7�t�� pu����� -��͏ۏ�����N� `�Ϗ��o����)�;� �����8���\�˟ ݟ����;�Q�گI����m��4�F�X��2TOLERENC�sB�	"�L��0�CS_CFG �( +x'dMC�:\��L%04dO.CSVY� cֿ�x#A ��CH�z _/x.�G��},���RC_OUT �)�- z/��SGN *��"��27-MAY�-25 14:3�8�����]� Z�t�����x.�����#�pa��m��PJP���k�VERSIO�N ��V�2.0.11~+E�FLOGIC 1�+� 	d���ٓ��p�PROG_ENB�2��WULS�' �p�_WRSTJN� ����p�MO_OPT_SL ?	��]�
 	R5�75x#?�74D�6E�7E�50i�d�o��2E�d��j�"�TO�  .����k�V�_� EX�d�%� �PATH A��A\��M�_�~+�ICT�F�,� '�`�e�g��}�STBF_TTS�(�	��Eмt`���0MAU�\�ߧ"MSW��- )���},t���.�! ��]l�R�v������4SBL_/FAULy�/��#>GPMSK�ߧ"/TDIA��0�����`���!12�34567890xS�l�P���� �//%/7/I/[/m/ /�/�/�/�/�/L0-PV �� �/�2?X?j?|?�? �?�?�?�?�?�?OO�0OBOTOfO8<x�UM�P$�I� �AT�R>�O�@PME����OY_TEMP��È�3��4���DUNI	�w�YN_BRK 1���x�EMGDI_S�TA	��_�LPNC�2_SCR 27[��_�_�_�_�& �_�_o o2or�nSUQ13y_+?|o�o�o�o�lRTd47[� Q��o�o���_>Pb t������� ��(�:�L�^�p��� ���� ?Ǐُ�0�,p ��+�=�O�a�s��� ������͟ߟ��� '�9�K�]�o������� ��ɯ�����#�5� G�Y�k�}�������ſ ׿�����1�C�U� g�yϋϝ�ׯ������ ��	��-�?�Q�c�u� �ߙ߽߫�������� �)�;�M�_�q��� �����������%� 7�I�[�m�������� ��������!3E W��{����� ��/ASe w������� //+/=/wa/s/�/ �/�/�/�/�/�/?? '?9?K?]?o?�?�?�? �?�?�?�?�?OK/5O GOYOkO}O�O�O�O�O �O�O�O__1_C_U_�g_y_�_�_�_�gETMODE 15'E�fa t�|�_GgRROR_PROG %�Z�%���HogTAB_LE  �[1O��o�o�o�ZRRSE�V_NUM �R?  ��Q�`�a_AUTO_ENB  u�SZdw_NO�a 6�[��Q�b  *�*6p�6p�6p�6p�`�+5pOastHI�S�cXa�P{_AL�M 17�[ �2��6|6`+t�@��&�8�J�x_�b.p  �[4q�R����PTCP_VE/R !�Z!6oZ��$EXTLOG_7REQ�v�y��SIZ�܄TOL�  XaDz�r��A ܄_BWD�o�%��fQ���_DIn?� 8'Et��TXa b[�STEP�g�y��P��OP_D�O�v$v`FEATURE 9'E�Q��QHa�ndlingTo�ol � DER� Engli�sh Dicti�onary�7 �(RAA V�is"� Mast�er���
TE�0�nalog I�/O��p1
�0�uto Sof�tware Upodateb� "/��k�matic B�ackup
�d�
!��gro�und Edit�B�  25LCameraT��FX� "Lo��e�llT��L, Pn��omm9�shۡ��h600��co�u���uct��p�p�ane� DIF����tyle s�electѡ- �/�Con��9�onOitor��Hd��tr�Relia�bT�ϣ(R-Diagnos���Q�	�H�Dual �Check Sa�fety UIF�c�Enhance�d Rob Se�rv��q �v�	ԸUser F�r���T_i�xt. DIO f��fi�� )�\�e�ndܰErru�L���  prנ*�r�O�� @���EN�FCTN Me�nuİv����.f}d`�TP In?�wfaco�  
E��G��p;�k Ex�cذg�C��Hi�gh-SpeܰS�ki��  Par�+�H���mmun�ic��ons��\ap��urf�?�X�?t\h8U��¯connZ�2Т �!�Incr��s�tr)�8��M-6��KAREL C�md. L��ua��}��B�Run-�Ti�Env�(P<�@�I�<�+��s���S/W�"H�License����� ad���ogB�ook(Sy>�m�)	���"MA�CROs,��/O/ffse\�f���бH�!�Y�M1�M�echStop �ProtZ�3� 5�
�Mi4�Shsif\��B6S�MixܰQ����H��Mode Swi7tchY�Mok����.�� ��Mt�Q�g��� �5��ult�i-T������)�P{osj�Regi>�^��  ! �PA��t Fun1��6�iB/��R�Num�Y�3�G�P/���� Adju��	�/g2HS�)� o(��8�tatu���A�D ��RDMޱo}t�scove&�� #e�v�㱗��u�est 867.��o�\���SNP�X b��Y���)�L�ibr%�
�rt �I���� "����.�S�o� ��s in� VCCM����� j�����㣀{/I�� 710�?TMILIBX�8���g�Acc�����C/2�TPTX<�� �Teln��Y�@����K�PC�Unexcept^ܰmotn�� ��������\m72�5����w�5��� � h640SP CSXC�i � j�*�� RIN��W9e���50,��svrl�زmen" ,��fiP-�a��㪼P��Grid{�play F O/�0�? ��ELR;�|�s20��ORDK��sciiw�loamd�41d�st��Patd��Cyc8T�h���oriɰ:ѽ7c Data� q	u6�2�0�*����܁��FRLam�c�K�HMI Deb��(����k�PC�����Passwor�d�644��Sp������D#YELLOW BO�	?1�wArc%�visu�4���#ti�Op�^��! 2��aO�pof�� t��ֶT1o�̸���HT��xy��	�   $�t�۠ig��10Ơ �41\+�JPN �ARCPSU PiR+�8b!OL0wSup�2fil� �!��E@-�;�cro�c�82��v���$ [12jSS0e4tex-� I�7�S�o��tf�ssag"�� e��У�P��,���� "Tc Vir�t��v�!����d�pn�
�J3�S�HADf0MOVE� T�MOS O� TԠget�_var fai�ls l�>PU~1E����� Hold �Bus %�h��V�IS UPDAT�E IRTORC�HMA A�{�vYWoELDTV S ]��DtS: R741��ouiPb}�y���BACKGROU�ND EDIT �"RC$REPTCD� CAN CRA�SH FRVR s62z1�SCra���s 2-D��r �) "��$FNO NOT RE���RED �` m ���JO� QUI�CKaPOP FL�EN m41S�L�oc��gRTIMQ�%�#�FPLN: \FG��pl m�r`��MD DEVIC�E ASSERT� WIT PCV�;PB�AN#aACC�ESS M .p�c��Jo��Qui�±�KbldmgU�SB$ ��t & _remov�� P�g�SMB NUL�� ;a|�FIX��C���ACHIN,QO�L�`MO OPT� ՠa��PPOSyT0�WDU C�nwQAdd�`ad��ք0io�2��$PZ�`W\0.$0`O��IN&�P:fix� CPMO-046 issueC��J/aO-�0�r13�0Т- ��vRSE�T VARIAB�LES-P{��R3D� m��view ed��M��&�ea����b��of FD��5P:N@x OSs-1y0`�h sc�ڎ�t��s t�lő�7 WA�PZ�3 ?CNT0 T�/�"�ImR�)�ca ��Pu��POT:W�henapewB�S�TY E�{1t��p�tKQdo GET�_�p �p��VMG�R LOl�REAd0C~QW�~1�(�l��s�gD�ECTpL�pING IMP�R�DR(p+PB�PR�OGRAM�ERI�PE:START=U� AIN-;�Ӡ}M/ASCIIzP�ÂOF Lq�DP�TTB: N�pML$me P���`�:x�mo&�all�W`!�ӤTorc�A��U�HC�iLpԸtuh�`n�@ ch��p/GEA�!�tou͐��RCal��k�S7ign`� ND�ԗ�Thresh12�3��`��09p : �MSG_P�+0e�r  �Q�Aܠz�eron��0 H385��RImA�n�[2D��rc�0I��gOMEa`�pONaP�5�  נSREG:FF-Д� ]�'���_KANJI��n���J��c�0asn d<�!OA immc ��INISITALIZATI����~1cwem����dr+�� LB A�UWqm�inim�rec�[�c!�R���m$�ro -1>ѮS�ܰAir��@ұJ�1pdET�w�� 5`?�I�ow� u��< se 1+lc��YbPM���p��Q���R`vR&�lu<\�3�Re 0�4q2�q1#���m <a��arn��ঁBo�x fo��*PRW�RI�PW�S��v�0�9 F�pup�d_e-rel2 d�p� j��`━bet{we��IND Q����igE sna�p|�us��spo� TME��TPD�#�DO�p#aHAN?DL 1\k�`vR��ȀD�ny�S�v��Yoperabiql� �T*�: H � l\p��Vq�b�R�R< p�a*�c&2O�`�FA,�.�-QV7.o f.v��GT��pi�s��� ɠt�mLine-R�emark �� �RM-�` W�#SP�ATH SA+PLOOS UIFc��+5f fig�pGLA����Vrp������=U�0ther�Vџ Trac���tW�\b�s7��d�t�4� n�@  ���3�:���dK�y��i�t k8�d�Pay�R![2]�ü1:� g��s��dow2�XQ��0IS�q�q�EMCHK EX�CE C���MF� +�Xah�� 3�5\k��)���QB�t���'b���[�c���e �`k�S�Џ BUGr��cD$`PETp���f��c4��0XPANS�I��DIG��@O�oPmetTCCRG� EN��CEME�NT�A M̀K �{�`H GUNC�HG �`� EXTЩP�2�bQS�93� wP8�x�ORYL�EAKq  H5�gyq�PLC WRoDN R �O /uN�QSPE=p��G*V ��$�tn72�0\3pGRI��A��rT�PMC E3TH��pSU7p�`�  j5/n�PE�NS�PN,��*P �ont�`BROW��`!sRMV AD�Dz CN qDC����PT3 ALA�2@ ���pSVGN? EARLY�R��ŰH57�GaJwLAYҀE (@MM�PPD�p*@H��S I`P�OUC�H8���V�F�q�c�omH�x ��ERR{OR� DE nJ���RO�CURS8pI��N4q��-158n7�RSR xP#aUp���Rqy�T�Fz�;�p0k��t�� gՂ��B�SY RUN�N�  a�`�BoRKCT�!RO�p�3@ \apSТ�A1XxP���h8+ q��ISSUr} sP\X�PTSI�K1�M10_�IPSA�FETY Ck�ECK[��Á����ഁ<#X�� �TWDp2�@�@�INV��OD ZOp�5X���t�DUALy� G"M6�0�"rF#��E��dPdNDE�X F�t*U�F�"Pʀ�0sFRVO117 A�PqT6�KtqFALP_TP2477D6_��P�!;HIG� CyC�t;SNPX� �MM��tq�d~�V�q�q#�
"��DE�TEC�Tq*@RR�U�qA�P�5p�9 By�)<9���7T�~�Pds� k��	���!Q���� t�\4A�;A0�2 "Ke@" 8@HI�qXF�8@4@H�PRDC"�
�aMB8@�IXF�b���zOX@8@���a�Gx}E�B�Ccscr�J�8@�NdctrldA.�A�NZE�A5��Q��!�`�Df8@�`m�W878�Q-;� ��/� rm`�
��PmR̠78�@RI8@0q�Q (~\Mp� �0t��!{B8@\tQ<OTX�St0�3hB3nO��Vtp�A�@LCF�L��� �Rplc�f���J8@�WTamaai�E8@mubov2_ miTA�O�S8@U`T[tT��AqPr674xSS�hape Gen(��8@j�I�[R�`�@b8@T����%q (u8@��II�^�Q~C�a��[8@;Ynrsg0�4�� � 4�CtMr68@�r5hB5�zVnr�etsp "r�P�o�wng0bGCR�E�Ka�ޠ�DA�T�E�k�crea#t.�q�M�a�oks>qgtpad1P��(�tputZj�{�������܆28@�����Q����sl�o��� �hexH�TB�88�ď�keyH�8@F�pmZb�NR�u7A+�nrgc8@UQ�pp�bUZ�dp0aj92�1xSpl.ColAlأcq�\A��RNq̩UA� (J�8@ip��_�WA��_�Y��a7�hB7�ͦtp[� "TCLS9oKb���clskyh[��s�pkckZd���$��TQ���dA�rx�71�0a- KAREL Use Sp�OFCTN9�a�7l�0s0a�� (���a��@~C8@��MI��c8hB8"   �8@� v	�v�	   lmatea99�qM��|��E�mcclm5�CLM;�� �j��E�3et���aLM	�h��yasp,���mc_mot�B�N��8@H����Q��su'��Q��p��䅮���joi#�xߕ��A_log�Z���trc�B����ve�ϓ�v��QWX��~6�finderxS�Center F81�lSw520��hal6rX� (<�r,�Q�Ձfi�Q �NH0�I�ۡ���A8@uL��t�q�a "FNDR�Vϳ���etguid�UID�C8@����������TA@�nuf;��P���ƞC�B��_z�Ӡo��qG��������l���fndrpTY��2䁴tcp"�,qCP MF�}3�8@517��6s38 �E��gf6��(���K��Q��-�X��A�t	m6�P�İ��Q���	�͘��t!m�Ĵ�b8@ej��TAiex��aP�Aa8�ذ�cprm�A�|�l�_vars� �
��dwc7 TS��/��6��ma7AF�Gr�oup| sk E?xchangJ 8@��VMASK H5~�0H593 H0a�H5@� 6� 58J�!9�!8\�!4�!	2���"(�/��;OPMI� `@a0hB0�0ՁU4U1#SK(x2H�Q�0I�h��)�mq��bWzR�Disp_layImQ@vJ�40�Q8aJ�!(P���;� 0a��0���� 40;�qvl "DQVL�D쌞�qvBXa`�uGHq�OsC>��avrdq�O��xEsim�K40sJst]��uDdX@TRgOyB�Bv40)�wA~����E�Easy No�rmal Uti�l(in�K�11 J553m�0b2v"�Q(lV40xU)���x�����k986#�8Uϕ�|�rP "NOR��dw d.a}oKksu�O�W���OY�W`��j0�6�H� menuuyP6�M�`wRX��R577V�90 ޛRJ989}�49�b\�`(�fity �����e�<?��Vsmh`��8��C0�Sv�q�8���w�pn "MHMN<� �ޣx�Ay`�o�3�u�`f�І�x�t��tRz`Q��LV��vP�tm��D�|I�1{oPx �2|�䎋I�3I/B�odstǏًmn����}/ensu_�L<����h!!��Rt��huserp��0Ҹ�ʐcM�_l�xP�oe����poper����xdetbo/�l>�x ���Ps$p�`���O~Pydspweb͓���z'R��u�Rr1C01&S՟{t�`2�Z4�30������`4�
�4�5��KQ�m8[T��dUCalG40 `�Q)p40}������9;��DA�� �v	LATAump�d�\bbk968&��68c�fbl�41969y�9�|�D����bd� "BBO�XêM��sche�d����m�setu0M:�����ff��� 40��n�41�ϒ�40q��col��|�1�xc�ؘ���li��X�0׀��j��&�8�4 <�r=o5�TP E�#6��ryK42r���;�(T+Q �Rec '�ʈ1Iw�84���ϼ�Ak971��7�1�;���parecjo��QNS�[T|���dXrail| nagek�M ,QT52 *� (���R%<x�80!bh�*��p��4��4�yDg�l�paxrmr "XRM�g�l�brf{���n��kl�~�9turbsp��p㧑- �l015	�g�625C�Mh�+ ���)89��	+��B�6��o�ҹ��x�7�q40����pd "TSPD�=��tsgl��l�:dQ0���8Bct���K�vrE�aܮ������  ��!���21�`( ?AAVM �2��0 �@fd TU�P him (�J545 l)��`8 616 %��VCAM ���CLIO (�0�:�5&  (F�\ MSC �Rt"P~BsSTYL��D!28 :2\ NRsE F2h SCH6�pDCSU �tpsh O�RSR �rD!04~�SEIOC& �\fxh 542 �LEX"� ESEaTn�8!H ��sh8 �7H �MAS�K�Ø"7>��OC%O*`x�!03"6�!�/400:66$ G63�9.6[8LCH!6O�PLGR703
5M'HCR��0C� (!� �06�A.f8!5q4
��00DSWb �588�180 �h!37 88 (D�"�02C24���27 	q9�25��2-6�0�5��9PRS�T bBFRD�MES�!zB�93�0 _ NBA � 6� HLB 3� (~!SM�@ C�on� SPVC ��8!20z��TC�P aram\?TMIL A��@�PACETPTX� �@p TELN� 96��29�%U�ECK��r UF�RM et�P!OsR ORP IPL%�CSXC�0j�1CVVF l FQHTTP stA"X)�I#� CGHP8Z?IGUI�0��hPPGS Tooml� H8�@djZ�0�!@�h!63�%�@532Q\�31 B�h!{96�%R651�R�s�!53 TFA�D�R41�8"1 V��oo�"9��41�775�"/@�P�VC�TO�@�U�!sh!8=0�%PRXY�R�!�770 �b8 88O5 ol3P� L� �аdi� �`ڳh L�CP{Q� TSS ��b�26:����@CP�E �HT@VRC8~�tQNL ��@�002 %��b	0d3is� �`7 <��a�\0�T�`1 �`en�b4 652�`)FU02Q0Πo`p�P�tu�r4 $r5�N��RU0p@nse��QJp1 APFI�[ Jp3�g34�g40 alxrE1t�44w46� ts U0  7v�0O��r�5�e�p7 p "�sw�a61:��r4,��r5 QpwGr`D�$�p8R�"sP`tQ�5b�36w77�w8`&�v83���r8�&:���pOq8�8 "rk�ey8�9F��a90�91 p�#@��� n�D095�g97*pur�A1@d���P�|P�q1�0QplSq1�p#4��]a!s1@s	l༂8�Ӽ�\1�d�1�`��v�@{�1t4p�ae��5 h2���`�6ޣ��7�f1 p@��d�YpCqd�ـd��1�`uq��� Cu1�< Oq� ��7ReU1$ �u1�Pϱ� ��@�- WQ158 �ase C��9 |B��60 82ń��p���4 (WaAi��`吢!��7E���8�EU1P`ro$9�<�1��<�2��<�@	0��T��l�5Jäl��cC���9%�M#CR��P�2�`�:Q2@967�Q��)8��9Z�2TPBh���P�2P7U5@�o���
�5�`U���3 w���?A�E�1��c�qAwl��A�|1��512 f��D1�u5Р���a5p�$��56�+a��Q5h��Ұ�1 @��ppz�b[�538 xa�B��|p�4�2�11�/q5�p�4U5�P16 (߲�Pz��0��8�P�����p�e�5`�e5(�/�P`b�bf>�X��$Z�U�5�d�\� X�7� 	  ��8 �k_kv��79 �s�82 &�H5@��E6���p����h���ñ���3J"�`���4 3Ȥ59ѧ6R�0t���8��6D0\$�$�4 7��!����<�j670\tchk<�Ps��<�B<�90��7�<���<�\K�<�q�Ӻ�A�C<���q�<���<�t6��sg<�lc���	FA<�H��<���<�����<�hk��<Щ� B<е�o�<���<��<K�<�dflr��<����� ��o�`���hD�;�<�gEvam����B<г�oќ����<а�KЀ�creexl����P��<��¬|���j6<�s��prs.`���\���<��7������fsgan��P�b�t�at���<�L��1B !�s�vsch/  �Se�rvo S��ul�e>�SVS��4�4�1u�_<��� (�����ched��,`��~��A\�� ��  B���B�qA�����cj�� � 5�1�<���Ә�p�css "ACS<�&(� �6� �����c �el���Q����t�orchms�<�- T�Ma`Ѵ����09 J5;59�8 J681s�7� 8��b��<Чa8����te,s������/�E�� m���ARC.�� �1q�4�!=��C�tc�pA�@t���f�S F����7#�2xуSE�r���Ut9mS�0960'����RC������� p��96G= '��"H5W����L���\f�� �PA Tb���`!4U�#!Stmt�E �0�� �pMA�!pp��z�2?�in_<�PX��r�X e/cW�����V����et�dl�vߏ\ove�to���܏��mmonitr�\���|#�0st��?.6a���PP���! pQ�!y`�`ame �ΘArol�c�43��0 �p���0�1� 25�  ��<� v	��v	�A@�818\n; <s�I�B|�2�pMPTP"�|�C�1mocol�� ,��CT�v�'!� �A��̴�8P53��y`Touchs�s�`��<��J5���Ѩ`mP����n[PQ�a,��E�a��IP&
�Pt	h�A<�KF#R�m;�Q�etth�THS�R'�q-�Rt��o "PGIO�#!$s�vISwka�"WK���!�MHqH54J��5w5n/�Sm/���@ 7�*�da��8�`!w/Ac��tsnf Tk�/�#gb�a��(u`��^m�`u��Z���ܱQp�є�#���HKa<��M��t5Q tZ�a<��dFS5GK�4���G�1or��dW��64��tPx���P ����x,��?$����P<�Z4e7�g �"SVGN.ox�copy "CO;��Wj$�O�A�9� "FSG�ѧ�%7��_��5f� wQSWF*!">(�sgatuɀ����_
��tp_TPiDo��9�79�#�dߎ?���h�GAT����!#��  �Гf�` ��"/� �w�Z� �b?6?� ��� �� ���E ���M� �chrT� �K6K� ��sms� �o6�ѐ�gtdmen?3 �?���� ���mkpdt�d2 ���, ���pd�Q�X� ����� ���m?vbkup. �[�xC�С��mkuno���prp���mklh �4��s �niU�<�� �ldvrw���glg�4�� ��棑���aut7�.p б�旐 �ַ������su3� �Ǜ� ��ȷ� ���\ �6�b2 X� ��&�� �����A�4�  ��B ?  946" ��f�B� �t\paic\p4k947 ����F#���� �ict3as���pa`���cc:�<��o�����'gen�� � ��F��lnp � ����st1f@��1��wbO�c��Ջ�`��߄�vri �ߢ�а�-T� ��<�p�flow� OP�Ac��ow���R�50qtS �#T� (A��4�#���pѣV�cu3�QF� ��SfI�ac����46�0���s&��pa��!!0���� ���55�b ��o)�p���0娿
�aOfcal3�P� ��f��}���`�f��m�	߳�p�d�m�/���a�/��$C`ѷ�� �!? track\P� �0�ine/Rai�l Tr�]TJ�699W�T  (L��8 (`љT.�`�%��D���P0� (��8�4A8��_ɛ�⇒4��P��� �3�b3����alV@ �NT`f���%��Iin]08m���aen���� ��&?5�c@Itst3@��$�� ��`�,R9�%���0��%��popen�ers-OW dD#ev��F�M�6W����|A�Pc"�l!es v� �,��R��V$�Q��0�U<�V$ �k9j ��6��# �����%pwaop/!OPNUp�V ��2celL��8g_��/�6��tscG��$��V!�3z� 5vrop����7`�n(`�V"2 D�a V'O$:S9��� PumpE��jQ��@�" ��!
��@бM SC#�@��)P��AC�`�x�� � v����� \mhplu�g�@g�"7P��uXK")㠱io7�CJ0���E�LIO q1�g 7A93շ�5� q9 t����4rb �ST��R��CPJ9s89�P�LSE�'� �e C3Q(P �/Ov���o�P� ?a I1�R���55���f�I1`�tcmio���MIO�����Ut}co1"CL01V� �cBK`io��uM?���Sl�I0�ߢ�DEg �o���f �tI4\onfdtI���ex%�p27�Inte�.TB CoMoo1E��R�(do554# (;r>Ex,��nR##ipc�/>��qp5���
oQé�1��p����7/o���ra�pd�CDV_��r�P�֮��qp2cnd(��s �p��a�o�r@`҄�S��"�c�a�c����2kIԿ?A�p�crt���or0�qd #��"���3p+���D�x�Џ��vr2k�0����AG�.+��c3ho�;�uC��(� �uV630�fwe  P�mී�@���`���TX�� ��d�ch�p "_��(	�3������8����\p3�v����ш�9�3��1 �����lo0w�[ͧ���chk���㳦s��s?Ө0�i�1h���2��i�w����s?1*�-	�:�O��vr������0�'���PFRAPW;at?1rneE�P�sp�& ac5� _A�rbo#�,�a��g@��������Qs<�ICSP+ 9_�x���� ��F��A9PH51IQ93 7��HX6hQ]PVR2`S5��fPR6 iQ�WPR� (P!am S�u�"�A�I>0�tpprg�0����`h�@2atk9�32�!��E�^��asc "8�C��S>i�atp�"�d�@1I��
g�dsblf�ltJA�Qsabl�e Fau�P{C�!��EV0ex/!DSOB (DC��t�$ �p��X 7� �� 5��Q�t3*�~���td9� "!%�(5��sb9኏���\	�6#���@5�p$D@�550-Adju�st PointO"tVJ�Rs�z�䐄���!�X_�Yj��0\sg��4��}7y��\ada�"AD�J���j�Qets{ha<�SHAP�sŭ'jpo�r4�t �!��$ ��C|�	T�k!bRPKAR�/Qiagnost�ì!O!vV66 �J`ew0�(�L���/�&krlde� ��PP���hU b$���r3�Pp?q��ODBG2C��� �@X�o�1U�� ���WT`�@ipJCM��aipper O�pv`1Se}78 (MH GF� ;" :�&##�� a�x�֕$��388C�����#��9.�9C��g##PPk�Q��8�!�_"$ �"��=0%�P��A $���_�#%0AQ�C~2 M�at.Handl�E��!= &�pq MPCLGET�0�1(�3 �Tt&P�Sٰ'�B�1� �B0����&p��H��PP  �'p��@�C7PP	 �TG�tD5�}m�q�Afhnd "F_R?  �����PP	   xT?Q��n�P(Pa��To�P����?�pmpaOx��JP ak925��!2`@O�JRpsQ`B�2�unLHP�Tgse�GSo1�O�W�Q�T��v !�R�Ptpx~���JRdmon.��@��V�!ns�hYvr�QJ�g�Q�o�jY��HS~7sl�f ��pen�PDnR(R&���ɐ823'��ٔq ���g� ���� 1�� St�� ? �c\sltQ �!|QE�P��a�rtPg��P�� �v��"SE�DG8�s0�qtdgY T����vP `ho�s`<`����qc�`g
�e` o�w�a�@o"�ile6�H�e �ȅnR�� �e! j517�>Ճ��J%��e�`��Q!4��Q&�L�!F��J�=�o�5�z/l1�7���_�œ��`C0~C�  ���LANG j��A��������gad���#�jp�.��4�Ē�ib���s�Ƒpa���&���?j539.f�,�Ru� EnvA
������3H�z�J9�����h�ФP
Ҕ���2�2����� (KL�n-TimФ�⠤��p��3�TS����\kl>�UTIL"o���~x�r "QMGl���!������1 "���S�T3�\kcmno��SФT2����ut�.�lreadc�}�exY�ܤ�r���\��l��Фw�30��2C�*� -�CӀD�E!Ĥ� .��C� �R CV̴�Ҁ�\p��Р���p�tb�ox��.�@�cyc�sL�:�RBTE�v�eriOPTANE���;ӕ�k�e��0��a�ߦ�hg�ߥ��DPN��gp.v���r�ptlit���0�4��te\�cy����tm�nu3`�r���5?UPDT��������駣��ite| �� swto�<,���oolB�F"��Y���Q��(q��gr3��䪒��"�䴁Aw������߳��s�������������l<S���bx "O�� ����l����P���A�l\t�� ���ø����	�Col�e!��R C��r���&r �m;`��Cha�ng�Lq�T1 �r�cm3�"��
� 6 ���"����sP7���"L��222���2D457x�� CCFM�|H��accda��Q�c' ��KÕ0���K!����mo!��� ,$Á��!"
��� �/�/����	Y�,$��)�,$sk����m rC%tS1,$+��k1�%unc.,$oñ��1��sub�������1��cce�5/!&@��-/?-W/i&vs� }/�%#�#�/�.C��/� C%
�@? U �&+���F:qt�
pDЃ{ D	  U��:7�Dxmov.��P��DPvc5Q�t�fr@PeC_UYge�obdtg_y[tu ���P���PTUt�P�S�x�_�^z�_�\va�r�_�\xy�_�[pcl`c�P���P�U�e�Pgripsuaoskuti���ovfinfpo}��o�jB�b�P���Qud\�a�X��Pc�\Rrp�Qn ƅ�P�v�P)tm#qƆ0�P�v�a+rog�a��p\Q�?a+rpal?a{�{spa���P�u�Q��t�_TZp�0�osip�kag3r�ovlclay(�:�t�pT�Ad�pu?a�c�A�������KtKa�P����q�Tf|rdm��{r#in#r���s� ��2���|s�Pd�v�t�v��v�h�0��ys�tn* џ�yt'�1��p��D�p�uϑ#�u!l�@o�W6�2�si�updl�]�o�vr�on��`1L�z�`\��r���il3$|l4��ǉ#q54FyB��Տg{�`���{wcmxס���wxfer�~UYtlk2pp߿�UYconv��siccnv�Qʯxag��H�Z�lct`ao�=�yp��׭nit0����3������  ��� v	�gv	$��alϑ#pm�r&�B�eWa� ��f�%������I�@�߬�u�ͬ�KamT�`f���c��w��roǁ@#�5�����?� sm� �y�a��y넑���� ��`����͐ϑ��p��m�Wa�1��� A�6�S�e�X��ψ�\Q }�����������ĥw� ��西߭���߮�#q 0��rs�ew���1��a��z긱n@�.�۲�;�d������ � � Ad	�T$�1 p! �P��e �e �	lf@C�@�s�/�  ?�����8� ��������reg.��C=��o99� ~@����$�FEAT_IND�EX  z �_�e� �ILECOMP �:���1!�!z$#SETUP2 ;1%�;"�  N� f!$#_AP2B�CK 1<1) � �)��/�/ # %�/�/e4 �/ �/>%�/$?�/H?�/U? ~??�?1?�?�?g?�? �? O2O�?VO�?zO�O O�O?O�OcO�O
_�O ._�OR_d_�O�__�_ �_M_�_q_oo�_<o �_`o�_mo�o%o�oIo �o�oo�o8J�o n�o��3�W� {�"��F��j�|� ���/�ď֏e����� �0���T��x���� ��=�ҟa������,� ��P�b�񟆯����� K��o�����:�ɯ ^�����#���G�ܿ �}�ϡ�6�H�׿lπ����ϝ���@)t P�x/ 2� *.cVR��߅�*��@߂�F�j�T��PC�rߛ߅�FR6:D����V���z�T  �!���K� ��q�S�*.Fߢ��	�Ӑ���^����STM ��'����S���iPe�ndant Pa'nelS���HI����9���U�������GIF0;��������JPG��;���]oR�
ARGNAME.DT�y�>�\"����Rc	PANE3L1Y�%>��e�w��2�A/� //���/�3_/�/@��/p/�/?�4�/�I?�7?�/?�?T�PEINS.XML�?>:\�?t?�1�Custom T?oolbar�?Q��PASSWOR�Dg?w�FRS:�\:O�? %Pa�ssword Config{OR��O SO�O�O��_�OB_T_ �Ox__�_�_=_�_a_ �_�_�_,o�_Po�_Io �oo�o9o�o�ooo �o(:�o^�o� #�G�k��� 6��Z�l������� ƏU��y������D� ӏh���a���-�Q� ��������@�R�� v����)�;�Я_��� ���*���N�ݯr��� ���7�̿޿m�ϑ� &ϵ�ǿ\�뿀��y� ��E���i���ߟ�4� ��X�j��ώ�߲�A� S���w����B��� f��ߊ��+���O��� ������>�����t� ���'�����]����� (��L��p� �5�Yk �$ �Z�~�� C�g�/�2/� V/���//�/?/�/ �/u/
?�/.?@?�/d? �/�?�?)?�?M?�?q? �?O�?<O�?5OrOO �O%O�O�O[O�OO_ &_�OJ_�On_�O_�_ 3_�_W_�_�_�_"o�_ FoXo�_|oo�o�o�`��$FILE_D�GBCK 1<����`��� ( �)
�SUMMARY.�DG�oblMD:��o*n`Dia�g Summar�y+8j
CONSLOG qn��=qConsol�e log�7k�pMEMCHEC�K��2��qM�emory Da�ta3�;g� {)}�HADOW(������C�Sha�dow Chan�ges���c-�?�)	FTP��蝏�=��qmme?nt TBD;�;g�0<�)ETHERNET0�`n�q�~���=qEthe�rnet �pfi�guration���B`%�DCSVR�F/��'�@�C�%�� verif�y allC��c1�p� �DIFF�8��0�ůD�%Z�diffǯ{��q��1������J� �X�q�|�	�CHGD�&�8�ͿD�!ܯ�����2Ŀ����R� `�yτ��GD�.�@���D�8����FY3�ϳ���Z� hρߌσGD$�6�H���D������UPDA�TES.$�
�ck�FRS:\"�c��>qUpdates� Listc�`{P�SRBWLD.C	M��blN��e��p�PS_ROBOWEL\�6o+�=�loa� �o����&���J���n� ����9��Jo�� �"��X�| #�G�k�d� 0�T���/� C/U/�y//�/�/>/ �/b/�/�/�/-?�/Q? �/b?�??�?:?�?�? p?O�?)O;O�?_O�? �OO|O�OHO�OlO�O _�O7_�O[_m_�O�_  _�_�_V_�_z_o�_ oEo�_io�_zo�o.o �oRo�o�o�o�oA S�ow�*�� `���+��O�� s������8�͏ߏn� ���'��� �]�쏁� �����F�۟j���� ��5�ğY�k������ ��B����x������C�үg�v��$FI�LE_N�PR]����Y�������MDON�LY 1<��U� 
 ��ۿ(� ��L��5���Y��}� ��ϳ�B�����x�� ��1�C���g��ϋ�� ����P���t�	��� ?���c�u���(�� ��^�������$�M� ��q� �����6���Z� ����%��I[����2����VISBCK����ų*.VD�*� �FR:\V�� Vision� VD file Vd������ �	/./�R/�v/�/ /�/;/�/_/q/?�/ *?<?�/`?�/�??�? �?I?�?m?OO�?8O �?\O�?�?�O!O�O�O �O�O{O_�O!_F_�O j_�O�_�_/_�_S_�_�w_�_o~�MR_G�RP 1=���LeC4  B�`	 ��lo~li`�۬B��D���fnӺ�MT� ��� ����e`i`a�o �khb�h�o�dcic�.M��2K���K% M��5�G�K�E���|�i`=��Lu?��>��[P;�/w?��Ӑ7�.l}>���>���>w����r����p=�l}F@ �qhq��y�~g�fF6��D�MqD��� BT��@����l}?pD��6����l���5�?�5��|�l}�B�H@B���B�u�B(g2�Bi��B=���l}Ae9�A��UB�\�A�G?A�BB̀l叐�A������A�܏e�P���t��
���A[@?A�@�IӘ��� �Ο��+��O�:��_���p�����eBH` �Ă���㟯��'�d�
��Z��WZ�Ôb/�FX
�A@����@�33@�N���\��[���ѿ��@��񿋯�*π�N�9�r�]ϖρ�<��G�=�<��m]<�+=~�m<c^���8eN7���7ѷ7�x7;��51�~���X�=�(�C2^`Yb`U�b`�����Fߪ`Үb` b`�0�����C�^o�߂o �o�߸o��o�� ]� (߁�l�������� ����#��G�2�k�V� {������������� ��1����-� )������� 0T?xc�� �����/')� '/M/_/q/8��/�// �/�/�/�/?#?
?G? 2?k?V?�?z?�?�?�? �?�?O�?1OOUO@O RO�OvO�O�O�O�O�� _��J����`_*�_ N�_�O�_�_�_�_o o'oMo8oqo\o�o�o �o�o�o�o�o�o7 "[Fjh�x �t��!��E�0� B�{�f�����Ï��� ҏ����A�,�e�,/ ���������/�J�� ��=�$�a�H�Z��� ������߯ʯ��� 9�$�]�H���l����� ɿ��ƿ���#��O�O V� _z�D_V_��z_�� �_���
�C�.�g� Rߋ�vߛ��߬����� 	���-��Q�<�N�� r��������� )��M�8�q�\����� ������������7 "[Fk�|�|� ���֟3�W Bg�t���� �/�///S/>/w/ b/�/�/�/�/�/�/�/ ??=?(?:?s?:�L� �?p��?�Ϧ� O��$O ��T?]OHOZO�O~O�O �O�O�O�O�O_5_ _ Y_D_}_h_�_�_�_�_ �_�_�_o��@o
�go *owo�o�o�o�o�o�o 	�o-*cN� r������� )�;�M������� ��ˏݏď��%�� I�4�F��j�����ǟ ���֟��!��E�0� i�T���x���ï�?�? ��O��?OO�t� >O������ѿ��ο� �+��O�:�s�^σ� �ϔ��ϸ������ � 9�$�6�o�6o��Zo�� R����������5� � Y�D�}�h������ �������
�C�U�� y�����d�����:��� ��+Q8u` ������� ;&_Jo�� ����//گ4/ ��x�j/4��/X�n/|� �/��/�/!??E?0? B?{?f?�?�?�?�?�? �?�?OOAO,OeOPO �OtO�O�O���O�O_ �O+__O_:___�_p_ �_�_�_�_�_�_o o oKo6oooZo�oZ��o �o�o�o��xo
G 2kR����� ����1��.�g� R���v�����ӏ��� 	��-��Q�/*/�� N/��r/�/ޟ�/��/ )�D�M�8�q�\����� �������گ���7� "�[�F�k���|����� ٿĿ���O�O�O��W� B�{�fϟϊ��Ϯ��� ������A�,�e�P� ��t߆߿ߪ��ߪo� �+�=�a��߅�p� ����������� � 9�$�]�H���l����� ����������#G�2W}h�p��$�FNO �������
F0� �  >#�1 D|�� �RM_CHKTY/P  � �q�� ��� ��OM�� _MIN� m�����  X�� SSB_CFG� >� ~�Jl�Aj�|�TP_DEF�_OW  m�|��IRCOM� ���$GENOV�RD_DO�ܠ��THR dz�d�_ENB�� �RAVC_?GRP 1?3� X�e/��/�/ �/�/�/�/�/�/? ? =?$?6?s?Z?�?~?�? �?�?�?�?O'OOKO 2OoO�OhO�O�O�O�O��O�O�ROU? E\� q���|���8�?#��O__K_m_o_ꐖ  D3���_E�_2q�@A��\Bȡ��Rp��>Y_6 SMT<#FC-�Ufoxo�o��HOSTC,1G�Y?��_ 	��h�k�o�f�oyeCUg y�z1�������p	anonymous�5�G�Y� k�w��o�o�o��� ���*�<��`�r� ������ˏ	���� �&�8����������� ���ȯگ���M�� 4�F�X�j�����ݟ�� Ŀֿ���I�[�m�� ��fϵ��ϜϮ����� }�����,�O�Pߟ� t߆ߘߪ߼���/� A�C�(�w�L�^�p�� ���ϸ���������� a�6�H�Z�l�~����� ������9� 2 DV��z���� ��#��
.@�� ������������ �//g</N/`/r/ �/����/�/�/? Qcu��/[?��? �?�?�?�?)/�?O"O 4OFOi?�/�/�O�O�O��O9m�aENT 1=H[ P!^O_  `_?_._ c_&_�_J_�_n_�_�_ �_o�_)o�_Mooqo 4o�oXojo�o�o�o�o �o7�om0� T�x����� 3��W��{�>���b� ��Տ���������A� �e�(�:���^������㟦�QUICCA0�̟ޟ?��1@��.����2��l�~��߯!ROUTE�R௼�ί/�!P�CJOG0��!�192.168�.0.10	��GN�AME !�J!?ROBOT���N�S_CFG 1G��I ��Auto-sta�rted/4FTP:?�Q?SOBχ? f�xϊϜϮ��?���� ���+�߿�P�b�t� �ߘ�6�����(� J� �1�C�U�g�6ߋ� ���������x�	�� -�?�Q�c� ?2?D?�� �������)�� M_q����:� ��%t����� m�������� ��!/3/E/W/z{/ /�/�/�/�/�/6H Z ?n/S?�w?�?�? �?�?�/�?�?OO<? =O�?aOsO�O�O�O�/ 
??.?0O_d?9_K_ ]_o_�_PO�_�_�_�_ �O�_�_#o5oGoYoko �O�O�O�O�_�o&_�o 1Cogy� ���oT��	�� -�|o�o�o�o����o ��Ϗ����)�;� M�_�q��������˟�ݟ�ÿT_ERR� I�����PDUSIZ  ^���$�>=�W�RD ?޵w���  guest+�}��������ůׯ��SCD_GROUP 2J�W �`�1���!��L_��� � ��!�	 i-y	�E���Q��E EATSWI�LIBk�+��ST� 4�@좰1��L�FRS�:аTTP_AU�TH 1K�<!�iPendan�������!KAREL:*���	�KC�.�@���VISION SET���u���!�ϣ��������	� �P�'�9߆�]�o޽�CTRL L���؃�
��?FFF9E3��u����DEFAUL�T��FANU�C Web Se/rver��
��e� w���j�|��������WR_CONF�IG MY��X����IDL_CPU_PC����B�x�6��BH�MIN'��;�?GNR_IO�K����"��NPT_S_IM_DOl�v��TPMODNTO�Ll� ��_PRT�Y��6��OLNK 1N�ذ��� 2DVh��MA�STEk�s�w�O>ñO_CFG��	�UO����CYC�LE���_AS�G 1O��ձ
 j+=Oas� ������//\r�NUMJ� �<J�� IPCH�x���RTRY_CN��n� ��SCRNO_UPDJ����$�1 �� �P�A���/���$J23_DSP_EN~���p�� OBPR�OC�#���	JOGv�1Q� @��d8�?� +�S? /?)3POSR�E?y�KANJI�_� Kl��3��#R������5�?�5CL�_LF�;"^/�0EY�LOGGIN� �q��K1$��$L�ANGUAGE YX�6�� vA��LG�"S�߀������x��i��@Z<𬄐'0u8������MC:\RSCH\00\���S@N_DISP T�t�w�K�I��gLOC��-�DzU��AzCOGBOOK U	L0��d���d�d��PXY�_�_ �_�_�_ nmh%i��	kU�Yr�Uho�zohS_BUFF [1V��|o2s� �o�R���oq��o�o# ,YPb��� �������(��U��D/0DCS }Xu] =���"l ao����ˏݏ�3n��IO 1Y	 �/,����,�<�N� `�t���������̟ޟ ���&�8�L�\�n����������ȯܯ�E�e�TM  [d �(�:�L�^�p����� ����ʿܿ� ��$� 6�H�Z�l�~ϐϢύdN�SEV� ]�TYP�$���)߄m�1RSK�!O�c>�"FL 1Z�� ����߯������ߘ��	�:�TP5@����A]NGNAMp�$�E��k�UPS P�GI|%�1�%x�_�LOAD0G �%Z%0_MO�V�e���MAXUALRM;'�I(��~���#� V�#a��CQ[x�8��n��"�t1060\	 �F�	�Ϣ����������� �� D'9ze ������� �R=va�� ������*// N/9/r/�/g/�/�/�/ �/�/?�/&??J?\? ??�?k?�?�?�?�?�? �?�?"O4OOXOCO|O _OqO�O�O�O�O�O_ �O0__T_7_I_�_u_ �_�_�_�_�_o�_,o���D_LDXDI�SAc���MEM�O_AP]�E ?=��
 �5i �o�o�o�o�o�o�o~��ISC 1]�� �oTd��\ no������ ���I�4�m��f� ��$���������!� �E�ƏT�f�:����� ß�����z��ܟA� ,�e�w�^������~� ����� �=���L� ^�2���������߿� r� �Կ9�$�]�o�(t�_MSTR ^��͂�SCD 1_xm�W���S������ �=�(�:�s�^ߗ߂� �ߦ�������� �9� $�]�H��l���� ��������#��G�2� W�}�h����������� ����
C.gR �v�����	 �-Q<u`r ������// '/M/8/q/\/�/�/�/��/�/s�MKCFG� `���/��L_TARM_2a��w2 �#�\`Y>G`METPU�T`�"����NDSP_CMNTs5p06�5�� b�΂�>�"1�?�4�5P�OSCF�7�>P�RPM�?�8PST�OL 1c2}4@p<#�
aA�!aE qOG]OO�O�O�O�O �O_�O�OA_#_5_w_ Y_k_�_�_�_�_�Q�1�SING_CHK�  +O$MODAQ73d
?�7:e�DEV 	��	�MC:MlHSI�ZEs0���eTA�SK %��%$�12345678�9 �o�egTRI�G 1e�� lf��%��?   0A$�ÜfYP�a,u���cEM_IN�F 1f>7� `)AT?&FV0E0N�}�)�qE0V1&�A3&B1&D2�&S0&C1S0}=�})ATZ�� �H�E��q9m��xAu���X�������� ������ v�)���я��П���� ���*��N����� 7�I�[�̯ן���9� &���\����g��� ��i�ڿ������ï4� �XϏ�iώ�A���m� ������߿�ѿB��� �ϊߜ�O������� �ߩ����>�%�b�t� 'ߘ�K�]�o߁���� �(�_�L���p�+����������.ONIT�OR�0G ?ak �  	EXESC1�#23E45�`789�#��x xx*x6x BxNxZxfxTrx22�2�U2�2�2�2�U2�2�2�3�3�3aR_G�RP_SV 1g��y�a(�Q��|;�?`f��97��?��?���@I�Hm�a_D�i�n�!PL_NA_ME !�5
 ��!Defau�lt Perso�nality (�from FD)� �$RR2� 1�h)deX)dh9�
!�1X d�/d/ v/�/�/�/�/�/�/�/ ??*?<?N?`?r?�? �?�?�?�?�82S/�? O O2ODOVOhOzO�O�Ob<�?�O�O�O�O _"_4_F_X_j_|_�_:LhR� 1m)9`{\b0 �_p�b�Q @D� M �Q?��S�Q?`��QaAI�Ez�  a@og;�	�l�R	 0D`4b@4c.a�P�Jd��Jd�Ki�K��J���J���J�4�J~��jEa�o-a�@���o�l�@�z��b�f�@�S���a�Q�o�c�=��N��
�����T;f��`���l��*  �_p  �$p> p��$p��o?p?�߆�������o�Bntr�Q`�skse�}�l�p��  �pu`oj  #p��v�ks�� 	'�� � �I�� �  ��ޮ}:�È6�È�=���N��b@^�d��n�Q���{�R��x���nN. �� � '���a�`@a�@�t�@p�@p@CpC�0�f0�+pB/pCz3}�P�@%��Ea�poo�$|m����gA%���. ���zc�u����QDe����˟��(��m��� �t O�� ru �4� �R�c��s�' :�u�a�P�`� �?�ff � �����7� ���گ쬛af��>搠���iP�P;�e��S�Ea4f�u�>L�X��s�b<	�I<�g�<#�
<�2��<D��<���
vo��¯�S���S.�c�?fff�?u�?&찗d@T����?�`?Uȩ?X�� ��Z���T:z�TB��W a�з*dů�ρϺϥ� �������&�8�#�\�h�+�F. Kߘ�G߀��3���Wɯ���G?�@ G���� X�C�|�g�y����� ����jZ���ￏQ� ���ߙ�����3��� ����/A��t�_������� ����F ��@+Fp�IP�t�e�%���[`B�0� ���<ze�cb�!@I�
�M`�B@��@`��9@y��?��h� �@�3��[N��N�N��E��<�/�:/L �>��ڟ��A�p�C��F@�S�b/DpX������@��t��%�h���`/qG��G�knF&�F׿�pE,8{�/ �F�ZG����F�nE��DE,ڏ�/� ����G��F7���F��ED��.��C?.?g?R?d? �?�?�?�?�?�?	O�? O?O*OcONO�OrO�O �O�O�O�O_�O)__ M_8_q_\_�_�_�_�_ �_�_�_o�_7o"o4o moXo�o|o�o�o�o�o �o�o3WB{ f������� ��A�,�Q�w�b��� �������Ώ��� =�(�a�L���p�����=(r!3�ji��r����ꕢ�3Ա�xڟ�y�4 ���<�y��P�2�D��&�jb^�p�1w?����������ʯ���ܯ� �s�P^�PD�c�`�m���@y�\������Ӱ�¿ Կ�����.�G� ���}ϳϡ���홍�@U�_�J���$�y.� @�v�d�z߈ߚ�x�4� �������� ��D�.��2� �$[�G�D[�^�B���B��CH� ^����q���@��������t�h�M�_�q�����������^�^�Y�m�2��
 ���� #5GYk}�������h*�� ���>�x}��$�MSKCFMAP�  ��� ����m�N"�ONREL  �6�9_�"EX_CFENBk
7�]�FNC�}JOGOVLIMk�duyd"KEY�k�"RUN���"SFSPDTYU��v_�SIGNk}T1�MOT�z"_�CE_GRP 1-n��9\���/ ���/�/4��/?�/2? �/'?h??�?C?�?�? y?�?�?�?O�?@ORO 	OvO-OoO�OcO�O�O �O_�O*_<_#_`_-��"TCOM_CF/G 1o/���_��_�_
|Q_ARC�_�6��UAP�_CPL�_�NO�CHECK ?/ 5�;h9o Ko]ooo�o�o�o�o�o �o�o�o#5GT�NO_WAIT_�LF'5y"NT�Q�p/���q_ER�R�!2q/_�� AR_���"�x:�L�dT_MO�s}r�}, �\?P_|��_�PARAM�rs/�������MW��� =e�345678901.� @�R�)�q���_������˟����ݛLW��3�E�؏i�cUM_?RSPACE,��������$ODRD�SP�SI&�OFF�SET_CART�oݨDIS�ݢPEN_FILE��I!�Q�v�POPTI�ON_IO���PWORK t�'� T�|�/�^�F� ��䖱Z���	 �m���A�����i�_DSBL  ��v���ޡRIENTTOj��C���8�ῠ�UT_SIM_D�J�6	��VàLCT u�}\���Q��W�_PEXE���RAT����� ���UP ve����������Ϭ*�8��$��2�#h�)deX)dh�>O�X dY�� �ߣߵ���������� !�3�E�W�i�{��� ����������2n�� )�;�M�_�q���������<����� +=Oas����X��� O��1m(?���(�.�g�}�"0 �д�u�  @D�  &�?��?р~H�D4  Ez�Z3;�	l	� 0ӀS@(SM� �i�i ��H)!H,��H8�Hm��G�	{G�8��6�MV��� �SC�)���)�����Ճ�*  �_p  � > �� ,�//)/ �B,�Btr�«{�H�¼�/���/�"�# �,�0 �� �  �� ߽pj  B ��&X�?MU	'� � 12�I� �  ����-=���8U?g;/�@}?�0 ~.ѱ�?;Ѳ���rH[N5��?  'M�XD�> C)�f)�J BN +��=%O7O�R��@D1�o�o$����JWAD0�J5�4�: �1�E &?�O�O#__G_2]��� �t �O� ru �4 ��R<�Uɳ� :�%Ё�р� �?�fAf��@[�_�_V_{��o~��18р"o0j>�P�Q6YPрZo�W�rAdS�%�>L�w0�#�<	�I<�g�<#�
<�2��<D��<��׍�l�_��ѳMb�@?fff�?�0?&p:T@T��q?�`?Uȩ?X�-q �iyBq5Ya ��gI�_���� ��!��E�W�B�{� ��d�����ՏLnp�Ώ/�ʈG�@ G��U�ȏy�d����� ��ӟ�������yB =� ��?p���/򏸯 �߯R���'�9��o N�`�����~�����ۿ
ƿ�B�ĮD�e��ֿ;�ҿ_�J�?�A�h�oϨϓϸ��D4	��b!�_@���� �ħ��Ŀ����%�@I��)�M`B@���@`�9@y���?�h	� ��@�3�[N���N�N�E���<�/Y�kЖ�>��ڟ�A��p�C�F@��S���pX������@�t���%�h��߉!G���GknF�&�FצpE�,8{�� F���ZG���F��nE�DE,�ڏ��ૐ�G���F7��F?��ED��Mf�� b�M��q������ �����(��8�^�I� ��m������������� ��$H3lW� {������ 2VAS�w� �����/.// R/=/v/a/�/�/�/�/ �/�/�/??<?'?`? K?p?�?�?�?�?�?�? O�?&OO#O\OGO�O�kO�O�O�O�N(]�3g�ji�O�a��	U�E3Ա��O_<q�4 ��%_7_<q��P�Q_c_ERj�b}_�_1w������]�Y�_�_oP�_1ol��P�bPcn~���o�O�o{_�o�oY�`��o�o, /;M#�f0o�� ���Y�et�~�i#�1�C�yM�_����� ������{bS�Ԏ���	�?�-�c�Mj2����$�VG�z}�Bh����B��CH� }�9�֟�����0�B���wl�~��������Ư�T����\��qQ��U
 ί�0�B�T�f�x� ��������ҿ����܇��� ��]{x}���$PARA�M_MENU ?�Յ� � DEF�PULSE�	�WAITTMOU�Tl�RCV� �SHELL_�WRK.$CUR�_STYLj�Ϋ�OPT����PT�B����C��R_DECSNw�Te'�!� 3�E�n�i�{ߍ߶߱� ����������F�A��USE_PROG %P�%B��V�CCR��UeXÚ��_HOST !FP�!�����Tt`���������4���_TIME�� �T��  A�GDEB�UG��P�V�GINP_FLMSK]���TR����PGAʹ� |�[���CH�����TYPEM�Y�A�;�Qzu� �����
 )RM_q��� ����/*/%/7/ I/r/m//�/�/�/�/��/?��WORD �?	��	RS���CPNS�E̺�>2JO���BT�E���TRACEgCTL�PՅZ�� {`" �a`{`�>q6DT� QxՅ�0�0�D��Sc�{a�0���2��Q�?�?�2�4D1�2#A�O.O�@ORFcA�bB`D	�`D
`D`D`D�`D`D`D`D
`D`D�9�O�O_ _,_>_P_b_t_�_�_ �_�_�_�_�_oo(o :oLo^opo�o�o�o�o �o�o�o $6H Zl~����� ��� �2�D�V�h� z�������ԏ��� 
��.�@�R�d�v��� ������П������9 �*�<�N�`�r����� ����̯ޯ���&� 8�J�\�n��������� ȿڿ����"�4�F� X�j�|ώϠϲ����� ������0�B�T�f� xߊߜ߮��������� ��,�>�P�b�t�� ������������ (�:�L�^�p������� �������� $6 �Fl~���� ��� 2DV hz������ �
//./@/R/d/v/ �/�/�/�/�/�/�/? ?*?<?N?`?r?�?�? �?�?�?�?�?OO&O 8OJO\OnO�O�O�O�O �O�O�O�O_"_4_F_ X_j_|_�_�_�_�_�_ �_�_oo0oBoTofo xoN�o�o�o�o�o�o ,>Pbt� �������� (�:�L�^�p������� ��ʏ܏� ��$�6� H�Z�l�~�������Ɵ ؟���� �2�D�V� h�z�������¯ԯ� ��
��.�@�R�d�v� ��������п���� �*�<�N�`�rτϖ���Ϻ����$PGT�RACELEN � ��  ��������_�UP y��e���������_CFG z���������<���Q�c�r�$�DEFSPD {/���������IN~'�TRL |/����8Lի�PE__CONFI+�}՟��<��x�LID(�~/�~�GRP 1���������@�
�=�[���A?�C�C
�XC)?��B��r������dL�z����~��� 	 r�8N�Oۤ� ´�����B������������A���> �6>�7�D_������� �='�=)�� ��������	B-���Q�M��� G Dz����
� �&L7p[� �����/��6/!/Z/��
V7�.10beta1�<�� B=q��"`ff@��"�>����!=�̽͏!A>ff�!@w�ff�"�\)�"D��?�  �!1@�!� �!Ap�#W��h/??*?<?K;�w����O/�?K/ �?�?�?�?O�?O>O )ObOMO�OqO�O�O�O �O�O_�O(__L_7_ p_[_m_�_�_�_��_  o�_$oo!oZoEo~o io�o�o�o�o�o�o�o� DQy{/�#F@ {yw}�y{ջy �-������/�Z? l?~?w���t�����я ���������O�:� s�^���������ߟ� ܟ� �9�$�]�H��� l�~����_ۯ��� ��5� �2�k�V���z� ����׿¿�����1� \n�j�|϶�� �����	�4�F�X�j� c�χߙ߄߽ߨ��� �����)��&�_�J� ��n��������� ��%��I�4�m�X��� ��ί����������! E0B{f�� ����H�Z� ��Vh�ϴϊ�� ��� �2�D�V�O/� s/^/�/�/�/�/�/�/ �/? ?9?$?6?o?Z? �?~?�?�?�?�?�?O �?5O OYODO}O�O�� �O�OtO�O�O_�O1_ _U_@_R_�_v_�_�_ �_�_�_"4FxBo |����o��o�o //0/B/;�__J �n������ �%��I�4�F��j� ����Ǐ���֏�!� �E�0�i��O^���N� ß՟�������A� ,�e�P�b��������� �o o2oTo.�hozo �o�����o��Ϳ�o
 گ'�֯K�6�o�Z� ��~Ϸ��ϴ������ ��5� �Y�D�Vߏ�z� �ߞ����������1� �Uy��:��� ������	���-��Q� <�u�`�r��������� ��T�f�x�n ��������� ���7"[Fj �������!/ /E/0/i/T/f/�/�/ �/�/�/�/?�//?A? l�e?w?&?�?�?�?�? �?�?�?OO=O(OaO LO�OpO�O�O����* �O_@RdZ_l_���$PLID_K�NOW_M  ~���A��TSV ��]�P�[? �_�_o�O&oo#o\o��B��SM_GRP� 1��Z� dI`~�oo$Cf~�d����D��TPbj�oLk�f�o "~�U�o>n2 T�~����� 7�4���p�D���R� ��ʏ����������6��
�T��*������QMR�c��mT�EGQK? GR��(�#��� [��/�A�S������� �����$����W�� +�=�O������������� ���S�Ͻ�S�T�a1 1��ڗ���P0� @����E�ϲ������ ���M�0�B�T�fߧ� �ߜ�����������7�P�,�m��2����N�A�<��z�3��������4���������5)�;�M�_���A6x���������7����������8(:�L��MAD  ����� ��PAR�NUM  ���Ko���SCH�
 ��
��S+UPD��xaq{��_CMP_�`� <P�z '�U�ER_wCHK����Z���RS���_�QG_MO� �%_�~�_RES_G����� ��v/{/�/ �/�/�/�/�/�/*?? N?A?r?e?w?J'��W,g/�?L%��?�?�? N#(��?OON#w�4O SOXON#��sO�O�ON#  �O�O�ON#d �O_<_N"V 1��Uua^�@cX��Pp�P_$@cW،P��P_@@cV��P�"THR_INR���pbA%d�VMASmS�_ Z�WMN�_��SMON_QUEUE ��e��`UȨ`�N�U�qN�V�2`END4a6/NiEXE]oNeW�BE\`>o/cOPT�IO;g?+2`PROGRAM %j�%1`O_�0bTA�SK_I��nOCFG �o�^9pDATAɓ�B{@ev2w��� ���z��+�=�O���s���������nzIWNFOɓ��}�!d r��!�3�E�W�i�{� ������ß՟���� �/�A�S�e�w�҇ބ���| �98q�DIT �Bׯj~WERFL~hwS~��RGADJ �^ƪA�  ,�?E��8��Q�IORIT�Y�W���MPD�SP�a�j�U�W�vT�OG��_TGp���Rj��TOE�P�1�ƫ (!�AF�PE5 ����!tcp��%��!ud�?�!�icm<�Q_��XYm_<q�Ƭ�Oq)� *������Op������������ <�#�5�r�Yߖ�}ߺ�@�߳������&�*�OPORT�a�Op�A%�_CAR�TREP~`Ʈ��S�KSTA�X!*SS�AV`�ƪ	2500H809u�PT毙䕣�ƫ�����`X#�$�6�^m�URGEU`B��6A)WFP�DO�V�2��W�q�?Q�WR�UP_DELAY� �Ưe�R_HOT�hwR%z�����R_NORMAL��n��6SEMI�:y�QSKI�P���X%�x 	������� �X%-;%[m E������ �!//E/W/i///y/ �/�/�/�/�/�/?�/ ?A?S?e?+?�?w?�? �?�?�?�?O�?+O=O�OO1U�$RBTI�F��NaRCVTM쒻���m@DCRڕ���AB�u�B��*A���j@`�!@��w{)�F����xA�/Ž������l�_� <	�I<�g�<#�
<2���<D��<��
+__{_�_)`�� �_�_�_�_�_ oo$o 6oHoZolo~oi_�o�o �o�o�o�o�o D V�_z����� ��
��.�@�R�= v�a����������� ׏�*�mN�`�r��� ������̟ޟ��� ��8�J�5�n�Y���}� ��ȯ�����A�"�4� F�X�j�|�������Ŀ ֿ�ӯ���0�B�-� f�Qϊ�m������� ����,�>�P�b�t� �ߘߪ߼ߧ������ ��(�:�%�^�A��� �ϸ������� ��$� 6�H�Z�l�~���{�� ���������� 2 Vh������ ��
.@R= O�s����� /�*/</`/r/�/ �/�/�/�/�/�/??�&?28�AGN_AT�C 1��K �AT&FV0�E02;ATD�P/6/9/2/�9p8ATA2>�,AT%G1�%B960k9W+++�?,�1H�?�,�AIO_TYPOE  EC/�4?REFPOS1� 1� K x	�O[H/O/�O �MNO`O�O�O�O_�O�C_�Og__d_�_+K2 1� KLON_�_�o�_*o�_5A3 1��_�_�_ o�o�o�o>@oS4 1�Woio�{o�o3W�oS5 1��o�oJ����jS6 1� ����]�H����S7 1��(�:��t��ݏ���S8 1�����Ϗ	���r����)�SMASK ;1� O  
���NɗXNO�?���1�.�8�1AMOTE � �.DN�_CFG� �U���5�0BP?L_RANGQ�K!�Y�POWER �Q5 a�SM_�DRYPRG �%�%R���ȥTA�RT ����U?ME_PROׯ��d�.D_EXEC_?ENB  �5]�GSPD=����Y3Θ�TDB����RM\ÿ��MT_ѐT���S�D0OBOT_NAME ��S�;9OB_OR�D_NUM ?���AH8�0�0I$�	���s	�\���ބ� ��e��	@̀}�D|��D0PC�_TIMEOUT��� xD0S232�n�1�Q; L�TEACH PENDAN��j�5���=Q�x0Ma�intenanc?e ConsK"-���"+�t4KCLS/C�}�6���|� No U�se�=[߹�F���N�PO�ќ�5�z_���CH_L@�3�U���	J��?MAVAIL`����+��]�I�SPAC�E1 2�=L ����p��扢�J@����8�?��� ���V�w� N�������������� �4�&G
l�}d	 Q5U1���������` 4&G
l}d(�#��2����� ���2A/b/%/ w/�//�/�3�� ��	/�/-/O/^??@B?�?�?�?�?�4�/ �/??&?�?J?l?{O��O_O�O�O�O�O�5 �?OO1OCO�OgO�O �_�_|_�_�_�_o�6_*_<_N_`_o�_ �_�o�o�o�o�o!�75oGoYoko}o+ �o�o����)��>��8Rdv�� H�����ӏ%�F�x-�[��G ��� R�;�
�� ����ԟ���
� �.�@����c���p���8�¯=�dؠ��ϟ ���!�3�E�W�i�_� q������x��կ� �'�9�K�]�oρ�w� �ϛ���Ͽѿ���� 5�G�Y�k�}ߏߡߗ���߻������ `S� @��8堯F�"�*ل����� �߇������,��� �V�h�2�<�N����� ��������.L 4v�R\n��Ĥ��
f�7�_M?ODE  ��M/S ���&�߂��Ïb��*	��&/�$CWORK�_AD]	1@,^�!R  ����t +/^ _INTV�AL]���hR_�OPTION�& �h�$SCAN_TIM\.�h��!R �(��30(�L8�����!��3���1�/@>.?���S22�41�9�d�4�1"3��@����?�?�?���IP���@���pJO\OnOE@D�� �O�O�O�O�O�O__�(_:_L_O���4X_�_�_��8�1��;�o�� 1���pc]�t���Di�1��  � lS2��15 17o Io[omoo�o�o�o�o �o�o�o!3EW i{����wc� ��	��-�?�Q�c� u���������Ϗ�� ��)�;�M�_��� `[����ğ֟���� �0�B�T�f�x����� ����ү�����$�7�  0��� om� �������ǿٿ��� �!�3�E�W�i�{ύ� �ϱ�������v��� /�A�S�e�w߉ߛ߭� ����������+�=� O�a�s�����ߖ� ���� ��$�6�H�Z� l�~������������� �� 2DVP�\�  �A����� ��%7I[ m�������/ �/C(/ N/`/r/�/�/�/�/�/�/�/?F;/?B?vF�x1 ;?�w=	12345�678{��l�@�P�?�?�?�?�?O9/2ODO VOhOzO�O�O�O�O�O �O-/
__._@_R_d_ v_�_�_�_�_�_�O�_ oo*o<oNo`oro�o �o�o�o�_�o�o &8J\n���o ������"�4� F�X�j�|������ď ֏�����0�B�T� f�����������ҟ� ����,�>�m�b�t� ��������ί����(��6yI�[�@��`���������Cz�  Bp*   ����254F��$�SCR_GRP �1�(�e@(�l��0�@ `1 �[1s	 )�3�C�<� t�vrY�8P�}�k�ܤ����95C����-u��ȡ����LR Mat�e 200iC Ə190�1Շ0LR2C �3�=OÆ��D�
f؜1u��2�U7��`1��v��@�u���	t�������h��$�^0�2� ��_2T�gϡϊ��o� F�D�f?��s���������ht ,Z���r�B�˰�P�N�g�rN�Aܰv�  @D���N�@����  ?� ��J�H˰��y�N�F@ F�`�� ����A,Qw b���n�N���`����B� �_J�n��� ��/�%//I/�΀E+:3��6?|?�5��
И/�/�#��@=�a��?��6B�07�590@7����EL_DEFAU�LT  I����� ^1M�IPOWERFL�  V�v5]2�0W7FDOk6 v5 ��ERVENT 1O���O�t3C��L!DUM_E�IP?�8�j!?AF_INEj0O��$!FT�?=N�OaO!Q�O ��PO�O!RPC_OMAIN�O�H��O��O�CVIS�O�I���OE_!TP8PP�U<_�9d4_�_!
�PMON_PROXY�_�6e�_�_XR�_�=f�_)o!R?DM_SRV*o�99gouo!RR8�o��4hdo�o!
�@M��_�<i�o!R�LSYNC4y�8�oY!ROS�?�|�4H�tO� 8c�����;�� _�&���J���n����� �ȏڏ7�I��m��4���X����7ICE�_KL ?%�;� (%SVCPRG1�����!�"�3*�/��4R�W�"�5z���6�����7ʯϯ�C��5�	9��oG�� ��o������D��� �l��񑔯�񑼯 7���_������ 4����]�������� ���'��տO���� w��%ϟ��M���� u����������?� A��Ͽ�ђ�؟ꐊ� ��ɱ��������?� *�c�N����������� ������);_ J�n����� �%I4mX �|�����/ �3//W/i/T/�/x/ �/�/�/�/�/�/?/?�?S?Ś_DEV ��9�MC�:[8�im4O�UT_Rf1~6i8REC 1���f0�0w f2	 [? �?�?OO;O&O_OmJ
 ����2W@�I�O �O�O�O�O�O�O_�O (_*_<_r_`_�_�_�_ �_�_�_�_oo$o&o 8onoPo~o�o�o�o�o �o�o"F4j Xz������ ���B�0�f�x�Z� �������������� ,��P�>�t�b����� ��Ο������(�� L�:�p���d�����ʯ ���ܯ��$�zO�Z� H�~�l�������ؿ�� ����2� �V�D�z� ��nϰϞ��������� ��.��>�d�R߈�v� �ߚ����������*� �:�`�N��f�x�� ���������&�8�� \�J�l�n��������� ������4"XF h�p����� �0B$fT��x�����5V �1��< PVOf1xQ�FO"!+f0f(}a?_TYPE�?�k2HELL_CFOG �z:f2/� Y+�/;8RSR�/�/�/?
?C?.? g?R?�?v?�?�?�?�?��?	O�?-O?OQN�/  �!%QOOP�O_B�L�A& �OL�B�@�#'gB2& �d�O�O�&HK 1��+ �OE_@_ R_d_�_�_�_�_�_�_ �_�_oo*o<oeo`o�ro�oa&�#OMM ���/�o�"FTOV_ENBr$!}*�OW_REG_U�I�oe"IMWAI�T�b�I${OUTrv$&yTIMuw��`VAL5>'s_UNIT�c�v�})MON_ALI�AS ?e�i ( he9���� &�8�&$�c�u����� D���Ϗ�����)� ;�M�_�q�������� ˟ݟ����%�7�� H�m������N�ǯٯ ������3�E�W�i� {�&�����ÿտ習� ��/�A��e�wω� �ϭ�X��������� ��=�O�a�s߅�0ߩ� �����ߊ����'�9� K���o�����b� �������#���G�Y� k�}���:��������� ��1CU y ����l��	 -�Qcu�2 ������/)/ ;/M/_/
/�/�/�/�/ �/v/�/??%?7?�/ [?m??�?<?�?�?�? �?�?�?!O3OEOWOiO O�O�O�O�O�O�O�O __/_�O@_e_w_�_ �_F_�_�_�_�_o�_ +o=oOoaosoo�o�o �o�o�o�o'9 �o]o���P�������s�$S�MON_DEFP�RO ����:� �*SYSTEM*  �l�*��RECALL ?�}:� ( �}�8copy vi�rt:\outp�ut\cal_t�cp.ls md�: over =�>1731461�12:15647�5 ����̏ޏ�t}1Bz�����tp~�������H�Z��;z�f�rs:orderfil.dat��tmpback\�=>laptop�-u9nqdge�h:12832 �6�ǟٟ�2��b:*.*��������>��P�b���6xz�:\ ����0�1�¯ԯg�7z�a��������C� U�h�z����0���ӿ ��������?�Q�c� v�	�Ϭ��������� �ϗ�*���M�_�r��� Ϩ�:������ϝ� &ϸ�I�[�nπ�ߤ� 6��������Ϗ�"ߴ��E�W�j�z���pr.pc��2�2�����h� zߌ��0�ASe�� �.���v�	� ���=Oa�� *�f�����( �K/]/p�/�8/ �/�/� �$�/G? Y?l~?�4?�?�? ��/�?�?COUOh/ z/O�/0O�O�O�O�/ �?�O.??_Q_c_v?_ _�?�_�_�_�?O�O *O�_Mo_orO�Oo�O :o�o�o�O�_�_&_�o I[n_�_�_6����tpdisc 0��c��=��O�a��tpconn 0 ��'� 9�ʏ܏��������H�Z��|�1��&� 8�ɟ۟� ������� G�Y�l�~��"�4�ů�ׯj}z���_dv.ls������C�U��_ �_o���o��ӿ�xo����o��?�Q�c�  ��$SNPX_A�SG 1�������� �P 0 '%�R[1]@1.Y1fϰ�?�p�%�� �Ͽ� �����6��@� l�Oߐ�s߅��ߩ��� ���� ���V�9�`� ��o���������� ���@�#�5�v�Y��� ������������ <`CU�y� �����&	0 \?�cu��� ��/�/F/)/P/ |/_/�/�/�/�/�/�/ ?�/0??%?f?I?p? �??�?�?�?�?�? O ,OOPO3OEO�OiO�O �O�O�O�O�O_�O _ L_/_p_S_e_�_�_�_ �_�_ o�_�_6oo@o loOo�oso�o�o�o�o �o�o V9` �o������ ��@�#�5�v�Y��� ����Џ��ŏ��� <��`�C�U���y��� ̟���ӟ�&�	�0� \�?���c�u������� �ϯ���F�)�P��|�_�x�PARAM� ����� ��	���P���p�OFT_K�B_CFG  �����״PIN_S_IM  ��̶��/�A�ϰx�RVQSTP_DSB��̲}Ϻ���SR ��	�� & ?CAL_DV�����ԶTOP_O�N_ERR  ������PTN �	��A���RING_PR�M�� ��VDT_GRP 1�����  	з��b� t߆ߘߪ߼������� �+�(�:�L�^�p�� ���������� �� $�6�H�Z�l�~����� ���������� 2 DV}z���� ���
C@R dv������ 	///*/</N/`/r/ �/�/�/�/�/�/�/? ?&?8?J?\?n?�?�? �?�?�?�?�?�?O"O 4O[OXOjO|O�O�O�O �O�O�O�O!__0_B_ T_f_x_�_�_�_�_�_ �_�_oo,o>oPobo to�o�o�o�o�o�o�o (:Lsp� ������ ���9�6�׳VPRG_�COUNT��8���d�ENB/�_��M��鴖�_UPD� 1�	�8  
M�������-�(� :�L�u�p��������� ʟܟ� ��$�M�H� Z�l���������ݯد ���%� �2�D�m�h� z�������¿Կ���� 
��E�@�R�dύψ� �Ϭ����������� *�<�e�`�r߄߭ߨ���������\�YSDOEBUGn�Ӏ� ��d��"�SP_PA�SSn�B?4�L�OG �΅ʹ� ���
�  ���� �
MC:�\`��a�_MPC f�΅����ҁ���� ҁ��SAV żi���� ����SV�TEM_TIME 1�΋ (�����������T1SVGUNYSɀo�'������ASK_OPTICONn�΅�������BCCFG ��΋O� H�2!`;A�I�r]o� ������8 J5nY�}�� ���/�4//X/@C/|/g/�/�/ ��, �/�/ ??�/�/H?3? l?W?�?��?��0�? �?�?O�?&OOJO8O ZO\OnO�O�O�O�O�O �O_�O _F_4_j_X_ �_|_�_�_�_�_�_o �X�  o2oPoboto�_ �o�o�o�o�o�o �o:(^L�p� ���� ��$�� H�6�X�~�l�����Ə ���؏�����D�2� h�o������ԟR� ����.��R�d�v� D����������Я� ���<�*�`�N���r� ������޿̿��&� �J�8�Z�\�nϤϒ� ��~������"�4߲� X�F�hߎ�|߲����� ��������B�0�R� T�f���������� ����>�,�b�P��� t������������� (��@Rp�� �����$6 ZH~l��� ���� //D/2/ h/V/x/�/�/�/�/�/ �/
?�/??.?d?R? �?>�?�?�?�?�?r? OO(ONO<OrO�O�O dO�O�O�O�O_�O_ _&_\_J_�_n_�_�_ �_�_�_�_�_"ooFo 4ojoXozo|o�o�o�o �o�? 0BT�o xf������ ���>�,�b�P�r� t���������Ώ�� (��8�^�L���p��� ��ʟ��ڟܟ�$�� H��o`�r�������2� دƯ����2��P���$TBCSG_�GRP 2����  ��P� 
 ?�  {���w�����տ���ѿ���/�A�T�[��~b�d0 �p�}?P�	 HBHA��L�͌�@�B   C���϶ˀ��ϟ�3D����A���x����A��T$�9��6Sff��f�@P�C��Ǝ�@�f߬��C� �ߐ߮ߴޥ���%�� %�D�W�"�4���j��|�������?Y������	V3.�00s�	lr2c��	*2�*�O��A� ��ѳ33P��d��� x�J�y� � ������T�JC�FG ���l� o������8�����= K
%�Kq\��� �����7" [Fj���� ���!//E/0/i/ T/f/�/�/�/�/�/�/ s���??(?�/[?F? k?�?|?�?�?�?�?�? O!O3O�?WOBO{OfO �O�OP�<��O��O�O �O0__T_B_x_f_�_ �_�_�_�_�_�_oo >o,oNoPobo�o�o�o �o�o�o�o:( ^L������h � ��$��H�6�l� Z�|�����Ə��֏؏ � ��D�V�h�z�4� ������ҟԟ�� 
�@�.�d�R���v��� �����Я���*�� :�<�N���r�����̿ ���޿ �&��>�P� b�ϒπϢϤ϶��� �����4�F�X�j�(� ��|߲ߠ�������� ���B�0�f�T��x� �����������,� �P�>�t�b������� ��������&( :p^����t� ����6$ZH ~l������ �/2/ /V/D/z/�/ �/�/j/�/�/�/�/? .??R?@?v?d?�?�? �?�?�?�?�?OO<O *O`ONOpO�O�O�O�O �O�O_�O__&_\_ �t_�_�_B_�_�_�_ �_�_"ooFo4ojo|o �o�o^o�o�o�o�o�o 0B�oxf� �������� >�,�b�P���t����� ����Ώ��(��L� :�\���p�����ʟ�� � ��_�*��_�l� Z���~�����į�د � �2���h�V��� z���¿Կ濠�
��� ��.�d�Rψ�vϬ� ���Ͼ������*�� N�<�r�`߂߄ߖ��� ��������8�&�H� n�\���>�����x� ������4�"�X�F�|� j��������������� 
Tfx�D ������ P>tb��� ����//:/(/ ^/L/n/p/�/�/�/�/ �/ ?�/$?6?��N?`? r??�?�?�?�?�?�? �? OODOVOhOzO8O��O�O�O�O�O�N  9PS V$_�R�$TBJOP_GRP 2��E��  G?�W<RCS�J\{��@0WP�R@T�P � �:�T�T �Q[R	 �BL  �U?Cр D*W[Q��_�_?fffe:�lB �P�f�f@`�33D  $a�U3o>g�_��_po�l�P�e9<�}bbY��?٪`�`$o�oUA��gD�`$�co�Qu>z9�P�Aa�P}@a���C�Z`xEp�o]A6ffpu�`aD/�U�h�� �r��~�a�RieAq�`�q��@9q�|�d�&`%���c333|D�\P8���?�`c?L�pAp[QB�b��k�}� ��z�� >��ffԁL��� T�f��fo ��Nw@� *�8�f���r�,���П ��ȟ��'����F�`�`J�X�����SC�V�ء��	V3.�00�Slr2c�T*��TQ��� E���E��A E��E���3E�iNE��!hE�فE�ۑ�E�I�E���E���E��rF�F��FM(F��5FBF�aOF�\F�"f,�z  E��@ E�� E��� E�  E}����� E���_�� EȆ�Ԏ��ᆰ� F  � F� F$� Fj` F�@� F�P F�`� 9�IR9�%o���L�_ �
�V��LQ��8TESTPARS��XUP9SHRk�A�BLE 1�J[$4�SV�+� �0�
V�V�V�WQV�	V�
V�Vȥ�QV�V�V�뱅�'RDI��TQ�϶� ��������f�On߀�@�ߜ߮����ކ�Sl�RS 0ړ������� �����#�5�G�Y�k� }�������������/] k�o��*	�%�7�I� ����+�=�O؆��NUM  �EUTQ�PP ��밆�_CFG �����Q@<PIM?EBF_TTq��8RS~�;VER�<zQ;R 1�J[O
 8�RP2� �@5  �� ����//&/8/ J/\/n/�/�/�/�/�/ �/#?�/?Y?4?F?\?Hj?|?{_�h@R�
<PMI_CHA�NG R �3DB'GLVQ`IR;Q��0ETHERADW ?�E;@�S ��?�?TO6V�0RO�UTe!JZ!��D�OwLSNMAS�K0HRSAA255�.�E��O�O8TOOLOFS_DIq���5IORQCTRL �s[���n]8]_�_�_�_�_�_ �_�_o"o4oFo�
�_�Tofo�og�PE_D�ETAIH3ZPON_SVOFF)_��cP_MON ��"P2�iSTRTCHK �J^�mO�bVTCOM�PAT�h;C�d�`FPROG %JZ�%CAL_DV� -=�m%QPLA�Yr��j_INST+_M�@ �|�g�t�USe]orLCK���{QUICKM�E�0)�orSCRE�F�3Jtps��or�a�f��2w��_{���ZyISR_�GRP 1�JY/ ؛ 6� ����;�)�_�M��8����Y������ �͕�����/��S� A�w�e�������ѯ�� �����=�+�M�s��	123456�78����f�X`�1��Ћ
 �}i�pnl/۰gen.htm������0�B�X�Pan�el setupF�}<�ϘϪϼ����� u�k��*�<� N�`�r��ϖ�ߺ��� ������ߝ�J�\� n�����I�?��� ���"�4�F���j��� ������������_�q� 0BTfx�� ����� >�bt����|3�~UALRM�p�G ?J[
  �*/!/R/E/v/ i/�/�/�/�/�/�/�/�??<?�SEV � �n6�E?CFG ��m�6���A�1   B��t
 =?�s3E�? �?�?OO+O=OOOaO�sO�O�Gz1ʂ��k� SΟ�OH7Isv?}{�`(%0?"_p_ I_4_m_X_�_|_�_�_ �_�_�_o�_3o�L�c �M�OAoI_E�HIST 1��i  ( k`���(/SOFT�PART/GEN�LINK?cur�rent=men�upage,153,1}o�o&�+�o�eedit��b�s�ou��(';�n2�o���*��5r�o�148,2�/�|��������S�,3���� �2���ӏ�b71쏁������� 6q)oߟ���'�9� ȟ]�o���������è�R��aR����%� 7�I�L�m�������� ǿV�����!�3�E� Կ�{ύϟϱ����� d�����/�A�S��� w߉ߛ߭߿���`�r� ��+�=�O�a��߅� ��������ʯܯ� '�9�K�]�o�r���� ��������|�#5 GYk}��� ����1CU gy����� �	/�-/?/Q/c/u/ �//�/�/�/�/�/? ���;?M?_?q?�?�? �/�?�?�?�?OO�? 7OIO[OmOO�O�O2O �O�O�O�O_!_�OE_ W_i_{_�_�_._�_�_ �_�_oo/o�_Soeo wo�o�o�o<o�o�o�o +?(?as� ����o���� '�9���o������� ��ɏX�����#�5� G�֏k�}�������ş T�f�����1�C�U� �y���������ӯb����	��-�?�Q�<���$UI_PAN�EDATA 1��������  	�}�/frh/cgt�p/wholed?ev.stmc����ӿ����)pri��.�Ip}2�V�h�0zόϞϰ� )���� �������0��T�;� xߊ�q߮ߕ���������Bv�� �   ��f@�E�W�i�{�� ������6������� /�A���e�w�^����� ����������+�O6s�l��  ��������� 1C�g���� ���L	///?/ &/c/u/\/�/�/�/�/ �/�/�/?�/;?M?� ��?�?�?�?�?�?0? Ot%O7OIO[OmOO �O�?�O�O�O�O�O_ �O3__W_i_P_�_t_ �_�_�_�_Z?l?o/o AoSoeowo�_�o�o O �o�o�o+�oO 6s�l���� ���'�9� �]�D� ���_o�oɏۏ��� �#�v�G��ok�}��� ����ş,������ �C�U�<�y�`����� ��ӯ����ޯ�-��� ��c�u���������� �T���)�;�M�_� q�ؿ��|ϹϠ����� �����7�I�0�m�T� �ߣߊ���:�L���� !�3�E�W��{�� � �����������r�/� �S�e�L���p����� ������ =$a����}�r�����)�*�� Vhz��� �����.//R/ 9/v/�/o/�/�/�/�/��/?�������$U�I_PANELI�NK 1����  � � ��}1234567890_? q?�?�?�?�?�4��]? �?�?OO1OCO�?gO�yO�O�O�O�OYIY0�:�M��[0-/S�OFTPART/�GENA1?CON�FIG=SING�LE&PRIM=�mainedit �OI_[_m_YJ_$_�M=wintpe�,1@_�_�_�_XK  �_$o6oHoZoloo o�o�o�o�o�o�o�o 
2DVhz� �������.� @�R�d�v��� ������Џ����M 0�,M9P E=Po�r?S�,Ico :�{�^�������˟ݟ �����7��[�m�P������O���BS0ߢ��C���/�%� 7�I�[�m�`C����� ��Ϳ߿񿀿�'�9� K�]�o��L���э͙� Q|����������!� ��;�M�_�q߃ߕߧ� 6���������%�� I�[�m����2��� �������!�3���W� i�{�������@����� ��/��Sew ����.���z� !E(W{^ ������/� //A/���͡Ϸ�}��� �/�/�/�/�/?�2? D?V?h?z?�??�?�? �?�?�?
OO�ϝϯ� dOvO�O�O�O�OE�O �O__*_<_N_�Or_ �_�_�_�_�_[_�_o o&o8oJo�_no�o�o �o�o�o�oio�o" 4FX�o|��� ��e���0�B� T�f����/������ ���ُ���>�P�3� t���i�����Ο��O/ �s/(��/L�^�p��� �������?ܯ� �� $�6�ůZ�l�~����� ��#O5OGO�� �2� D�V�h���Ϟϰ��� ����u�
��.�@�R� d�v�ߚ߬߾����� �߃��*�<�N�`�r� ����������� ��&�8�J�\�n���� ������������m�" 4ßXjM�q� �����B T7x������ A��//,/>/P/C� t/�/�/�/�/�/�/o/ ??(?:?L?^?Ϳ߿ �?�?�?�?�? OO �?6OHOZOlO~O�OO �O�O�O�O�O_�O2_ D_V_h_z_�_�_-_�_ �_�_�_
oo�_@oRo dovo�o�o)o�o�o�o �o*�oN`r �����m� �&�8��\�n�Q��� u���ȏ������"���?�?�{��$U�I_POSTYP�E  �5/� 	k�{���_QUICKMEN  ��j������RESTORE �1ו5  ��/
�2�D�h�mc�������¯ ԯw���
��.�@�� d�v�������W���˿ ݿO��*�<�N�`�� �ϖϨϺ����ρ�� �&�8�J���W�i�{� �϶��������ߡ�"� 4�F�X�j����� ����ߋ����y�+� T�f�x�����?����� ������,>Pb t������ (�L^p� ��I��� //ވ�SCREܐ?��u1sc�-�u2M$3M$4�M$5M$6M$7M$8<M!��USER/ 4/2F"T. O#ksW#�$U4�$5�$6�$7�$�8�!��NDO_C�FG ؜�  �,� ��PDAT�E �)��None V��S�EUFRAME � 
��&,1RTOL_ABRT7?���N3ENBX?I8G�RP 1�!��?Cz  A��3�1���?�?�?�?�?FO"OG:ېUx81g;?MSK  {5�A�g;N41%a��B%���O��VISCA�ND_MAXyE�I�c8�@FAILO_IMGy@f����#�8�@IMREG�NUMyG
�KRS�IZyC,���$�,SONTMOU4W0{D�%�VU�#_�c�� �P�2�FR:\�O �� MC:�\XS\LOG�VB@4 !�O�_�Q��_o
�z �MCV�_�SUDM10fEX9k
�f�TwV�2ۜ��p(��o=��͓o��j �o�o�o�o�o�o�o  2DVhz��K_PO64_?S�0Π�n6�uQ0LI� Q�z�x�qV� �|�f@�w�� =	��xSZV�~�����wWAI��DST�AT ܛ;�@�_ď֏�$����E�P12DWP  ��P G/����q��AP-��B_JMP�ERR 1ݜ�
�  � 2345678901����� ��ʟ��ϟ��$�� H�;�l�_�q����LT@MLOW���P�@�Pg_TI_X�('�@�MPHASE  �53��CSH�IFTUB1~k
 <���Ob��A� g���w���ֿ����� ����T�+�=ϊ�a� s��ϗϩ�������π>��'�t�K�!��#���:	VSFT1֣sV�@M�� ��5��4 �0��UA_�  B8����E��0p�����Ҫ�ӌe@��ME*�{D�'����q��&%�!�M��$�~k��9@�$�~�TDINENDcXdHz�Ox@[O��aZ®�S����yE����G����2�����������REL�E�y?w�^_pVz�_ACTIV���H��0A ��K��B�#&��RD�p��
1Y?BOX ��-�V���2�D��190.0.�� 83��254��2�p��&��r�obot�ԟ   pN g�pc� �{��v�x���$%ZA+BC�3�=,{� 낆;-!/^/E/W/i/ {/�/�/�/�/�/?�/ 6??/?l?!ZAT����