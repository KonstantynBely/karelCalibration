��  L��A��*SYST�EM*��V7.7�0107 10�/3/2018 A]  �����ABSPOS�_GRP_T �   $PA�RAM  �  �ALRM_RECOV1�   $AL]MOENB��]�ONiI M_IF�1 D $ENABLE k �LAST_^  �d�U�K}M�AX� $LDE�BUG@  
�GPCOUPLE�D1 $[PP�_PROCES0S � �1���UREQ1 � $SOFT; �T_ID�TOT�AL_EQ� $�,NO/PS_�SPI_INDE���$DX�SC�REEN_NAM�E �SI�GNj��&P�K_FI� 	�$THKY�PA�NE7  	$DUMMY12� ��3�4�GR�G_STR1 � $TIT�/$I��1&��$�$�$5&6�&7&8&9'0 ''�%!'�%5'�1?'1I' &]'2�h"H SBN_C�FG1  8 �$CNV_JN�T_* �DATA�_CMNT�!$�FLAGSL*C�HECK��AT�_CELLSETUP  P� HOME_IO�� %:3MACR=OF2REPRO8�/DRUNCD�i2�SMp5H UTOB�ACKU0� �	DEVIC�#TIh�$D�FD�ST�0B� 3$INTERV�AL�DISP_�UNIT��0_D�O�6ERR�9FR�_Fa�ING�RES�!Y0Q_<�3t4C_WA�4�1^2JOFF_� N�3wDEL_HLOG�28�jA�2?�1k@ơ?�� �����MOTOR_CEO 	 h Y0M_Ct� � 	�BREV�DgBIL�GGXI0~�BR 
 [ �OD<0�A	$NO� Ms0�@�DR2�!YW �V�AQ�B_D�# �d $CARD�_E�@T�$FSSB_TYPi�� CHKBD_S�E�5AGN G�� $SLOT_'NUMZ�QP�A�C��G �1_EDI}T1 � h1�G=H0S?@f%�$EPY$O�Pc iAP_O�KsRUS�P_CRrQ$�4�VAZ0/LACIwY1Db��Pk �1COMME>c@$D@fVa@`� ���QL*;OU�R ,�@�1HV1AB0~ OLx�ePz CAM_;�1 xCQg$�ATTR��P0A�NN�P�IMG_�HEIGHrQsWoIDTH�VTC�Re�0F_ASP�ECrQ$M@E�XP;$� Fv��CF\T X '$GR� � S!1Np=B_@NFLI<pwt
UIREs3��Q�OMqWITCH�vsQpN.0SXt�cG�0 � 
$WARNM'@f��P�� LI? �qNST�� CORN��1F�LTR�uTRAT�@0T�pAP$AC�C�1�  �� �OcRId`|S�{RTq0�_SF� ,�WCHGI1R�Tspu3II�TYJ�2 q�K*2 �`��p� 1sR*HD��cJ* �ȁ2Æ3�Æ4Æ5Æ6Æ7�Æ8Æ9���O�$ <� l~�xh�s1�`OIT_ 2�  4� ST�Y�w2Ge!VAR��)Y0���P��p��$ ��P��2�@�2�0+P��0'`?�yOJu4TOCO�3{PE�USH_��CE�p������EX�T9�E�a�E� 1 2 
o�.� ə 2P�����2@0��  H ip�Q�@1𕃗�p�4O O��q_�s�0o�� ~�ʘ
:�b�M<�r��g��@n�TWRIGz�dP���@0��j@A��5�P��6���w!�_MO�Rx� tW�FL�Ev�NG�1pTBA� .s㴴Q꺸�߸VP�BQ��P`�0�p�A0�v�p`�P�2� W�%��J%�_R�k�hPr�QJ(�vȑ�J��D�C���}�w�ul����P_}0OF� �  @� RO�����PqIT8C�NOM	_�0�1"�q3W ���$ �4����x1P٥}E�RAG�0�� �0��	�?R
$T�F����MD3�TD�&@U=0��Pb�YH�2{�T1��E,�� �u��v��v����PDBG4q� U��`PU�����4���:�AXc��rbET;AI�3BUFnV��)��!  |�p9��p[PI�b�P��EM��M��+���F��SIMQS����h�a�����MCµ1!~��@~0JB�pL�}1D�A���@� �%���" � �PN�S_EMP��$G�Є��P_��q3��1_FP:���TC ��9p�r��q0�s������� V�QAR�!h����JR!0ARSEGF�RA'�v 0qR�T�_LIN�S$PV!F�����,�#2R��D��a*)B��F�$( '�Ϝv�u�c ӳ�a=�.0m��M��	=�SIZ$� ���T����

�aRSINFz����) �p@��<
 <�� Lh�8�Ў�qCRC�uFCCC�pr
 ���} ��LrA���q��]"�D�t�s�C�j@�֐��$ pP�ٰ+(E�V+&�zFA!_��FR��Nm&����bі��#A1���!%c ��@s߻RGG`D��)�F �b��D<�24�LEW �As}�Ұ�ߒ.!�R_t&x 3�E������҃QR���`Ch�$LG�p���1Z`ѰlP�BPqA?@ٰ.�Z�R�"���3P�s�3)�8RA���3AZ���8' ��Od�FC�bApQp�F�p�4�)�s�ADILKWqOE�0/r�0ٱ@�p>D�p�p.s��S�P�x�0q�QMP.�`Y�C��0���U�baU���'��TIT�!��S��%V�n��D�BPXWO^��(��$SKdюR"�wDBTf0TRL��)˲A&`���0�`���DJ�ā�_CAL`�QbWPh@_WPLnLaߒD�a|W�a|W�Mh�DB�1��*Rv��PRc 
#P8��v���+ �����$��$� �L�Y,�_�S���q-�_d� .o�dENE��!/�;o�S�P�ORb0�H b�On 7+$L�c,$�S���0�k+ ��ձO�0_9DwA��ROS�r�� [�d�Z��cN�G��e�PA+�[�/ETU�RN�b�MRt�A�TU�pB�CR:�E�WM��GNA9L���$LA��Mu�;�-$Pj�.3$P@��/ap�Qb�C|t-ӶDO7 �j��d�a��fGO_3AW����MO�pڭB#PCS��1<mQISZ0�@֣��@���r5�qDᣐ��r������q��qW���NTV���rVE}���w�f�փ���Jm&�����SAF�E9ա�_SV�BEOXCLU�����"'ONL��ȃY_�yz��En4HI_Vv@>�PPLY_�m�VRFY_[S���r<r@��_ 2a`Px��w��� ��SGz  3R�
$$�*pGq�� X�;����B���V[�u�l�A�NNUN碓��I%D��U�bŃTp� �����b@��Ֆ"QE�F�pI5b4�$1F���D�OTJp�a� $DUMMAY�Q��� �#P|m0�u5 ` �HE�6U��W�уRr�k SUFFI	�A�pZP�!nP"�5��6��RMSW�u6{ 8�KEYI�-TM�a�ӡ,qΦIN<�հ"Qr@�t�7 D��HOST�P!��P���0 �����EM����k��PSBL� UL�R8 S�6z�=��PT|`Ʊ9 � �$���uSAMP�Z Ս��D��O I��`H�L�$SUB ����4`�]ၲ�C��SAV������ �3�s@�܀��P$`E�<APYN_B
S:� 0�DI��nPO�U�F��C$��R_�I; �ENC'2_S�0P;Qs@�����¸@Ń@��Ä-pQ<R�����a|����=  ��z���`pK�ddAn���AVERˡ���(Δ�DSP���PC�8۪�B/�Uѣ���V7ALU�HE@��MX�IP����OP5P~0 .�TH���#D��}�SY@-Ս�F;����d��w��@.SC�8����ET�$�>��FULL_DU����Dp����1g�Ư�OT�B�q�`NO�AUTOQ?	�!$R�S���Q�C��a�C>R/0�C1O�L @H *a�L�@�#� ����$�`������ ��Q��<��校�櫡���7��8��9��0T����1��1��1�U1�1�1)�16��1C�2Q�2����2���2�2�2�2�)�26�2C�3Q�3R��3����3�3�U3�3)�36�3C��4Q���SE�RA� <11�'S��Â1I`��^�v��FDӐ��B L�V1�!�V2]� igN�-REG&��GqE.p8pPC ,_��? �p�0?Q�к�E�p��B���"PD?��$TPA$VA�RIg��UP2f*�E 0���TD�� ��#x��,'&%!Q��wBACRF T����D)�L���P� IFI��P� �@<0*~%P;B��F)p��>PGt ;���2�� ST���!�@a� �`�&�/0	�"C+4	7P���s1�%�1(� 47FO�RCEUPl���F�LUS�H�Bp�_�E�2�D_CM�pE��h45IN_pY3m�^�
8REM]FŁ71�5�P62�0�8��:K�9Nw��8EF1Fӿ4�pINC�62wOVMIOVAI�TROV<N17DT<�HDTMXkL�0 H�pkJ҆P�H�5�C,�P62CL0_���Jȱ`k��9_Q��8_T�k0�KQ��pAL�Dz@42 X���Q�6�F�Xa`RQ44^IT�_�-�#0M"E��C9L��ıRIV���nREAR�IO�5#PC���@7B�r
8cCMJp0� dA�GCLF+S�QDY��X�@ב�S5T�ED�G01"E`e��FS9S�P�H P�=a�a����_<aSh<a�1��E�c<a3uk5�uf�GRAE �$I� ���W�ON<��cBEBUGp��b��4��p��_E �J ���H��T�ERM�eK�e[��'ORI�1�`Lv��GSM_ꀹ��`Mw/ �TA,yN�e���UP��O� -�q��Ju��csp�K$SEGxz	`E�L��USE�pNFI�!�r��a%�t�otL$UF}�H�C$U����p(�A��w�`T��� �NST�pPAT��a��PTHJ��&���V �r5���up��J��q�RELN�-�SHF�T�Ңq�@�_SH�OR	�#�+v 6p$�Ew��N1� OVRHj�-���Iq�qTU�= �AYLO��RC�I�R[����h��ERV��݁0��� �w�pN�w� 8��� �R�QPi�ASYMu�i�qWJ�w�&PAE�<�h��)�U��@�pB�@�p�(�V�Ph�X��hл�OR�pM�#��`SMT�%P�`�GR5 �c�PA��p���� �Q �� �(r!TOC�q�P��� $O�P�"(���
� �DQOR1ӰRE_�R��s-����� ef�R����z�X�x$e$P�WRZPIM���R�_U�{���r R�bHi% �_ADD�RH_LENG����
�M�R00S.H�S HS��;��wI��I���I��S�E[An��S3�#�T $��M�~1_OsFF[Ґ�PRMU�� N!HTT�P_T�H��U (��OBJ�R�x$-$LE�ĳ���V � ��AKB_!QT��S�lq3� LV��KR�R���H���BG>�LO0��	Q��p�Q2�w��'x�SS@��HQW=�q��WD����INCPU�bVISIO��-�����_����m���� �IO�LNZ"X�UPC^b1$SL���0oPUT_Z�$���P�P"���~0F_�ASCbY` $L u �u!���0U+p����q��e��߀HY`��fӡ�A�UOm0BcZ `RЫ��B }Ԋ@���ѧ�Pq3�����ф�������UeJ�&[�!NE���JOG�w,�DIS�2��K��	0Bc\ �Q��qV�j�CTyRR�j�FLAG�bv� LGAd] �0P��ҶcLG_SIZ�5 �� ��I���FD��I������ �� p���q���9��  9�I�9���9� p9�z@SCH_/ �Ŋ��SLNK��^��v1AERb!��� U�����L���DAU��EA����A������GHB���U�BOO>Z"_h Al�� �IT+�`h�REC1
SCR�0<�m��DIg�S�p00RG �"�Qh5�`�`��W�U�S��T�WoU����`�JGM�MNC�H�#U�FNKEY��K�PRG�	UqF����FWD��HL3STP�
V`��p�# �RSkHԐ]�C��I��`ӃP��U��� �����u�G�	i�CPO'N^IM��FOCU(RGE]X\�TUI�I��{"��#��#� ���A�P�R�N��8O�1�$ANAUқr�sPVAIL�CL��Ql�DCS_HI�d2_�2O8�Q4�S=P/58S+8�I�GN�� �����Tva�+
_BU@�@�`e�ĀT�"$��FP���r���A��ae�Ā��è���p" 1�52�53��1�7"0@�b � ����u(�B(ԓID_@�P؂��O�@C�qNFST��R���Y&p��q@ a$EFCK���ĎF�FEA�@�c L��{߰`�؎�X�g�����j���駨O_ d ����c�O0S�`C��e =�@CLDP��l�TRQLI ��:�dYRTFLGzBRP�aĆS�!DY�W��LD8�UpT�UORG:� �R����X_��m�BT�df ��`pT�aTJ�US�TdP�`�`��P?djaJcRCLMCUd�_�_gi��Ga�a9It��g d��"A�RQ�c$DSTB�:�E@ �f�hA�Xl� �h�lEXGCES�rbM��JhP�bl��eԳ�@�i���f_A@�j��X{�o�h�`K���j \��GROUܿ���$MB��LI�ܱ�sREQUIR��ro��|O�{DEB�U"�aL�@M\�k@
�J���sUb�a#ND��,�@�l����o�B�DCI"��IN�ʰ������L�\�W0N�8bq���`,�PS�TD� m��LOC%FRI��%E��%E�A"�&A�a�aODA�Q\�n X��ON��F����	�KI�B�U�U/������1FX�`IGG/ o �`�Cq�<��C��DR0�%oCk����{��Њ�wpu�DAT	A�7ǐE����0q����N�2p t W$MD�Iݱ)��C0��a��H؀$� �x����ANSW`�P�g�W!�D��)䂸�=`@�q +pC�U��V?��P��RR2�r Dհ�.��ADa d$CA�LI�`R�G�!��2N��RIN��<��'NTE
��2sy�楰8����
�_Nt@�����d�Dru�7DIV�fDHp�:ve�$V��[�vEA$�$Zӂ��Q�0ӂ�����w�H �$BEL�Tn��AACCEL�C1����ŰIRC��Ѐ�Ф�TcA���$PSpWRL   %���lS�۷��� ܶPATH��1�ѳ1�3 �q_�1��b��h�Bb�0C���_M=G�$DD��ܰ_$FW��ڐ�����ѳ����DE��P�PABN�ROTSPEEx��1��"`�J���1D��`�� ��$USE_���#P����SY����Ba �r�YN�`A O�OsFF�O�MOU��3NG�"�OL!�|�INC^�Ձ�¥��bx�׀`�bENCS������b�����d��IN�WBI ���@�b�V�E�Ы��23_UyPy��LOWL71A�C�"`��3�D�@�b�p� P��erC�����MOSd0|tMO���/pBgPERCH  P�OVG�KҒ� %A��pA6�dpAۃ�� �`�p;�?�40Ve�Wp���L�$��yw�����UP����1�L�TR�K��SBAYLOA 1Q��Tqa� �p�e�րd@��RTIXq��d@MO�����bTr�P~��d�ç�|�3��2���DUM2\�S_BCKLSH_C � ��r�q��WӉ����
fѨ�aCLAL��0��+a��#@NCH�K"`[ESx�RTY@L�#�ӭ5�Qّ_jCNf�_UMXp�	C�Γ�SCL���LM?T_J1_L�P�`�(��E�� �p� ���SPC0k���9��PC����!HP�p�šCc`RsXT����CN_¢N���ѳSx0F���V9�ZC�շ�m ��2qC�0�SHjC¢ �����Q���֣�d���>%���PA���_	P���_eP� h���0"ax�${JGw2}$�!�OG���TORQU+�ON^����`�r|������"_W��a�_q�5w�5}�5UI;I#;I}�F�� 1J�ab8a��VC"��0�d�b�21�>p8�?�b�5JRK�<�2��6=`DBL_SMt��;bMY�_DLw�;bGRV4Dw�D}��1H_P#�34�;J�COSHK��HHLN �0kK�5rDw�mI}�mI ?1�J�L]1�5Zf@|���1MYtA�HTBTH|ZMYTHET0<�NK23}�2Rq�u@[CB7VCBq�C�a�r\R?4jQw�jQ7VSqBw��RBUGTS4q��C�!Ձ?#�DV �Tx�C�W�C$DUx  yx�Q�����b�V���a9Q��ۆ$NE1t@�AIv@��b�U$�$U�&QA*USe\g:EEHEA�LPHXu1b�1bS �5�c�E�c�E1b�F�c(�j�FU�VuhVjhg���lV�jV�kV�kV��kV�kV�kV�iH�uh�f�r�m!�x�kH��kH�kH�kH�kH*�iOflOuhO ��nUO�jO�kO�kO�kUO�kO�kO�FF1b�WQ���E��hgSPBALANCE_�A��LE�PH_*US�P롈F��F��FPFULC�6��6��E��1s��UTOy_s �%T1T2w���2NZ�����&�@��8�`²���T"��OK�ı� INSE9G��U�REV��U����DIFK��1tl�I�1u>�OB��>CǩMI�e�4?LCHWAR�²��ABZ!��$ME�CH`Q�@�t��AXn�P��LgX�l��v 
���!����ROB��CR �Х���+�MSK_|�x P ��_)�R��x���M�1�������V�INݑ�MT�COM_Ct0��y�  ��
����$NORE��i���F�X�z 8� GRl�"y�SD(`ABz��$XYZ_DAxia���DEBUݑX}�F���{ �$G�wCOD- Բ���z���$BU�FINDX� � ıMOR��| $a�Uɱ]���v���7�G��} �� $SIMU�L� ۰���T���O�BJE�T�ADJ�USr�e�AY_I��!��D�ǻ��w�_[FIz�=�T�  ���ǯ�*���������p��DD�FRI4���T
RO� ���E1-�6�OPWO��0��~0�SY�SBU�`��$SO!PL��SW�UV���PRUNH�}�PA��D|�x�Q���_O�U�1q�*���$^��IMAG-���`P�IM/���I�N�0����RGOVCRD��n�]���P�����)`L_j�� �L��RB�*`2�M!?�ED�z� J"NC�M^�!�����SL��� x $OVSL��wSDI*�DEX�@����m1����V0��N���!�����������M!A �7� �_�SET� ��� @0� �RIV� 
�_dQ �9�,�6���p�� � Hx��y�z ATUS��$TRC`����Nt�BTM}�g�I�х��4 S�\���� D��E�Л�q�Lp�E�r��: > r�EXEx��D������b	�� �w�UP�����$+���XNN���m1��|1�� �P�GV���1UB�f�6�f�:�JMP�WAI�P��~L�O� ��F�S�$�RCVFAIL_C����R�������}� �Ű��@R_{PL:�DBTB�!����BWD�q�UM� �IG���Н�� TNL�� R��^�E��H���ODEFSP�� �� L����g_8jx�xUNI�Ӣ��v#R����@_L*�Pp�t�PI����а� v����ర��:�N'�KET�����P��� h~��ARSIZEE М ����!Sp�OR~:�FORMATc��
COz�!ߒEM2��4$�UX;������PLI��� � $S�P_SWIG����0� ~AL_ ��JuA-�BB�\PC-��D��$E���� C_9� �� � (5-��!J�3�P-�+�TIA4��)5�)6-�MOM�)�	3)33)3#3S�B� AD	3M63M6#3PUkPNR.4z53�z5#2ay!���?� A$PI(f�% ��$D�5!C�5.C�5 mT�6�;�T�T��V���ܡ����SPEED�pG�"ZD�g aFg�� ��aF�CpHp�I��SAM�����DaG�C�MOV ��TQ���UTeQg1;�/T2;�%�*Ґ0U� ��H��SINb\� �CiX�[`T��kZ�X�T�[�[GAM�M߆a��$GE�T����|�D�$0�
���LIBR7I.��$HI _�р�$�@fE� MhAGnj`[fLWBm�flji�f�[f�"��H��A� $PDCK;�D��|�_�@'�0�^R �)�!QUw)3tM6y~�# �$I8�R��D.�V�!�X�LE8��@�x�(Yp�u%4��0�P~ґUR_SCR)��q��C�S_SAV�E_D%��uNO� C@��$�pd�* �6�O��9���H�8� ��.�'Fu�EP�!���@ b�U8W$R<�[HQ� kF�HهՅ��Qt6�x M�5� �! �QW���2s*����p����W
�'�T�J� `�~0H�r�MŰx��CLw�w M�qC � $PY� �@�$W��[�NG ���!���$���$���$ ���$� +�=�#`�#|�J� X�O�#�!Z+�8w ���� p��S�3s�6�/�A�S�e�t@��!_Y�� |�� �)�p)9�3�#3�p�:���:E��e �޿ģ�r���t� ŤP$!�PM���QU�@ � 8��QCOU5q��Q�THƠHOL��Q7HYS; ESQ���UEw��r�OT��  �Pd�8e@�U�Ny�z� O O�°0� P��ִ�8�q��7ROG?���
;�2��O �յ��#�޹�INFO?ѕ �ư�I�:��u!O�IL (KpSLEQRFt�FEt��汒�D� �0����`O��`PSC?aE}`N9U�Ǿ�AUT�q��COPYQ �̯��M��N�����C��>� �RGAD�J��"XS���$�W�8�W�WU�P�U؍pW�jCG�kEX�� YCӒ�!D�NS�S� �$ALG�O�c��NYQ_FREQ��W�PEF��I$>�LAus��S�$3�PSECRE ��A�IF���NA�A%&�_Gusk�Q�˸ATf� ���*�R���P��mr�4���EL}Er  � ��!�NABӒ� EASI��قRN���SA�q��NP*`I-�t��`iq��� �s�ABx�� E�n@VXp-�B�AS�"/�*buTRp�� �Q��$F�n�c�c��ip���ߛ X �� 2��U�T��x���D�w��������'OTO�W�M ǰ_B�!��
�	)�>�ԝ � &�� p��3�64SRVF�1)S��C T_Om �\�3�	��5*�	6�	7�	8k�ѹS�r�0� @�M�C_F��<!��L�q�q�Y�R��� hP��3P���� ,KpFLА�q�pSYN� MM��C��PWRU�P��0=�ĲDELA�F�Y� AD���  ��QSKIP�5� i�C װO��NT'Q��P_װ ���p ����.C�;C��  �� �� �� �� ��� �9hq�J2�R^@�0� 4��EX`T�ӎ!=�ˁ�!���R�!'�R��RD]C��� ���R_�ORv�FUpQ�*���">�TRGEAR�亃�mrFLGl��ƠE�R��C<ç�UM�_� {�J2TH2�N�3" 1� ��!G��T�` I�R�w0M^1]�I\�D�REFQ1�q� lQ��1��_1ΐTPEbp��EG�� ���1��S�2ݳNbP5��2�О42�2��?@�?�?�?�?OG3�2�)O;OMO_OqO�OG4�2��O�O�O�O�O _G5�2�#_5_G_PY_k_}_G6�2��_@�_�_�_�_�_G7�2�o/oAoSoeowoG8�2��o�o�o�o�oL�oESMu�̠�n0�3��3E�qR�EMOO༴�� `��r��ˁ�sIO.Ѣ�yIUpˀ��R@W;ER�� _�L��!�s̠�G�$�DSB��A�9�W�R�TzC^0ˀ�RS�232�u���T�D?EVICEUH�̈́>ʂPARIT��W�OPBIT����CONTRްˁ�1���ʂCU����U�Xs�s��0ERFA�Cr�Z�[�I�CH�Ѳ L�������C��EFRO�M��{�GET_@� k�����pTu��ȔJ�PӀ�ѳ�� !x$USA@P|�(y�Ы�4�O����R8႒,�_O�NP{�����WR�K;M|�ὗ��SvF�RIENDF����$UF�����TO�OL�MY��$�LENGTH_VT�FIR��+����~�E@�9�UFIN�V*� �qRGyI��v�AITI�b2�X�A���G2���G1�0~�����P�����O_p��������$�C��	�TCp?�A�ȡ��G*0Z��д� s�p� 󪞘W��W�Ѥ�p|��E��X ]�*��L��T��H( �� �О�p�C�R�W����	��ɴD���`�`��ٱ��$�B��p���0��1ʘ���2��2-�3��3 ʚ�t�˙;ɐ�Sv�И\���h�$V� @�V��V� @� ������ چÌpb� �� ����c��V���pV�?��1au$A� �D�PR� E�[���S�!v�)!F�D��ҷ 0Io���� �ķ�A�pC���0�
�սS�q� ���R�Y����$RUNMN�pAX���A��L&����THIC²�K�:��1FE�REN����IF_CH����I��E�Sv��G1`�d�Rpk������_JF��PR\����RV|�A��ѹ2}�2 �VA�L�  ���� ���r��  2� ��S� U��d� �$E0�5L2G�ROU�q�TOT����DSP,�JO1G�񖂷 _P���AO�� A�ĆK4��_MIR��j�ȠML����AP��`EP08���M1SYS�s�vM1PG��BRK�(�,�,�Icqp��0�������ADՁ��BSOC ��pN�DUMMY14����SV��DE_�OP��SFSPD�_OVR/�C�� WZ�ORe5pN�k�fF,�fE�OV�H�SF�
�О^�F��t�l�̣��s�L�CH}�RECOQVV��E�W�ME �H�RO��(T�_����� @22s�VsER���OFSs�C��w�WD	{�(h���B TR��|�q��E_FDO���MB_CM�q�B8�BL��h���rԁV ���&�-В3�G���AM�����0/_M���)0�s�=8$CA;�)0D:��B HBK*��W!IO��f%�q�PPAZ*�!k)�$~%�%�r=DVC_DBv��!:�%�� t�"�%1�*0#�%3�&6ATIOs��2s�VqU��:��vCABQ� ��ѣ��G��E��_���SUBCP	U$�R�SՐ����+�\��7��� ���$HW_C#@�����7�A����l$U�NIT��l�1AT�TRI<��2R�CY{CL�NECA,2���FLTR_2_�FI]�9�23+�L�P^�=�<�_SCT6��F_�7F_�<B�JFS*���2CH�AՑgG�A����BRSD:&�	�%��p;_T�PRO0����EMkp_%��8�B�� �B��3U�DI`��RAIL�AC�#7�M��LO �4��(�661Ѭ650#PR� S���ОQC�!e�	/F�UNC��>�RIN�%�-���HP�T��RA�PA� B �S�P$��SWAR|�C BL ��WdAkAhh�DA���QRhceL�D�J �zc���Q(�zcTI0Қe���;$v�RIA��t�+AF�0P|��c(��e:�߲�#NCMOI�0�DF_$��'���LM�FA�HwRDY��ORG`�H�@����Z`uMU�LSE$� �7��G ��RT���p�$�$��$�� ����U��7� x��EG���J �qAR'�;320�9���u>`��AXE./�ROB,�W~���_�}SY���q��:�S$�WRI��|91;�0STR+�����q E�1��M�zS����Bq�<x���2 � OT}��P	$(ARY,�hQ4���]�FI��s�$�LINKq�ρ���_n�<L�y���XYZZ! ����'OFFD΂���%��B*�RT�P�PU�FI@n���0MB�TE�_JW���8oۃ�OP_����5����TB��Wrݒ�CB@��DUZK�6{UTURN��0��`���Q��H"ŗFL��@� K3�p4��t�7<^R 1���KQ�	M�K�8{U�50Қ7lORQV�Q�Sv� �s)���x�
p1��Us:7�T��OVE ��Ms@w�}s��s��r�W�M1��0��� �PsA�`����Y��" w�������s��>���QERV��Q	REA���S�A����r���UR��YaV6YaAX ��Ya5Ѿ�9���9� ��9ǀ�F�֐F��F� n�Fʔ�F��pF�S�F� pC�pS�pc�ps� p��p��p��p���p������DEBU�3$�Q�a1T��Y0򂏗�P�PABYWW! ����HP��
���# ��մ1�����-��� ֑�����n��ה�����q�d���bЂU�LABk�ť�0�#�:�� �+�SE�RVENB� �� $0��PA�!��POKO �����	��_MRA � d ��Ee�EcRRC;C�`TY�@�%�IJ Vk�5��TOQ4�r�L�p5�@����p���q �� p��T����E0_�V1��7�_�;Sl�2Be�2t���x������~#$W$@����i_������$�@R�`5���?�Z	�pFZN_CFG�p� 4�0w��@���3'�x� �` �>���s� � ���@	$2q���@`�FA�`���fdXE�D�`	/��q���0�PM2�pHEL�L��� 5�n0B_BASY3R�SR���P�sS��1�a� 1��%�2�3456�78�ROaO�`Հ��NL�q��AB��QP� AC-K��IN��Tr@i1�萾�Pp�A�_PUfYCCO�p��OU��P
`
aP�@BU7�TPFWD_KA1R�� ��RE��/pqP0`aPQUE��P�B@L4CSTOPI_AL������^S��3����SEMȤ3�$�3M�@� TYf�SO� TtDI��
@"`!U7�a_TM>�3MANRQ�&���Ec@Ss$KEY?SWITCH^SAA��!L4HEB@BEAiT"QQE�pLE
�TI8U#F�$"T@�%�O_HOM�`On�SREF�PR�QP&��^��Cc0OyC�`ECO�ි�`�`�IOCM�p'�!��p@��� DH��2 U��^"M�bx4"��FORC#fc =��OM�p � @���c�@Ud�P�p1eF�T�p�3eF4��NPX_�AS�� 0 A�DD2 4$SI}Z!$VAR.MpTIP��Cj@AKB���S���@�2$�P�rS"�qC�VOFRIF%���SH ZI�4�@NF�"�p� n��� x��SI#��TEO�Ԣn�SGL`QT݂@�&$0yS��<,�aPSTMTM��S�P�pD�BW�bTS�HOW�U&��SV|p�t�� ���A00>�ٱ�Rn@�W@x@�W�@�W�@�W5�YU6�Y7�Y8�Y9�YA�Y�p�WY@�W_��V{��WF�XS��h�Y�� �hi,��h)i��hCi����h]i1ji1wi1��i1�i1�i1�i2��Y2�Y2i2i2�i2)i26i2Ci2�Pi2]i2ji2wi2��i2�i2�i2�i3��y3�Y3i3i3�i3)i36i3Ci3�Pi3]i3ji3wi3��i3�i3�i3�i4��y4�Y4i4i4�i4)i46i4Ci4�Pi4]i4ji4wi4��i4�i4�i4�i5��y5�Y5i5i5�i5)i56i5Ci5�Pi5]i5ji5wi5��i5�i5�i5�i6��y6�Y6i6i6�i6)i66i6Ci6�Pi6]i6ji6wi6��i6�i6�i6�i7��y7�Y7i7i7�i7)i76i7Ci7�Pi7]i7ji7wi7*d�7�i7~�7�d��VPG0UPD��ˏ  @�0
�?�YSLO�� � �E� ��4W�G�}0հv0����AL1U��&CU����=F��ID_L�#���HI��I9B$FI�LE_�"�$$�3��SA��� h���N�E_BLCK�K#[�{Qd�D_CPUtٳ@t٧@%�7�x��T0�R �P�g
PWOP� ��LA/2S��������RUN~��������0~�"���"��� ��TBC�CE��X -$I�LEN@�#V�#I����I�!� LOW_AXI�K#F1I��2��M����|BP�I� 9,��TORQ!I�"��D���?PLu �2��I���[0_MA��@������TCV�>���T�!?�^�T�@���������J���M���J'�P��)����U�2�/0�������q JK��V�K�!�!3��J�0
JJJJAAL
@ @ �:4V5|^�N1�e�q 0���L��_��Q@��0E��� =`X�GROU��|Q��"BG@NFLIC��C� REQUIRE�4EBUy3E���@D�2��AF��DἛ@�S� \�;A�PPR� C�G�
vD EN?CLO�OS_MCP� d��y
D��E� �3@�MC�^���_M	G9A�C�POгq0��BRK�NO�L� ��PR� _L!I�1���J �PB������^���g��6/%nQ2"8���!�� ��p�]��'j�#PATH�'�!�#�!u�h�#�@Ұ�CNu0�CAB�@�INFH�UC����0C��UM8Y���C2���E]�3:j�3: �@P�AYLOA�J2=Lk�R_AN(�t3�L��~9z1n9�1�R_F2LSHR&A�4LO41�73�7>3ACRL_�A5��07f4��H��E��$H�&BFLEX�BC�JH�� :U�g���WGnDj�`����s���F1nA �E�G��������� � RE
��.�@�R�d� v������X�T�������@h������mA��T5g�QX�0����CT}X ���e~X	-? C L:^gy��
AB>�� � �����l�AT�F���CELWP{ �t�J� ��JE�CTR,1�ATNPF�v�HAND_VB�RqBA���$� $I`�F2�nX ��SW�)�`r��� '$$M�0�R�h�@�x��Pk�"��A�� k0������A���
�A�A�����Ъ�D�D�P� G��T�ST�\��\�N�DY�=��� ƅ|00�7nA�7�1m7 ��+d�@x`�P7%@% I%R%[%d%m%v#AC�$� ^�CD�"}�Y�<q��ASYM�%�P	� �&װ��-�1�/_SH�7 4
-��@/�*?<?N?`?r3Jy<�* �:J�@��9�D_V�I���q��V_�UNI�3���c�1J ��Ų�Ų�<ɴ�5ִ ���=���9* OOMŒ�c3D;C�`q$H���1�(�{�ENL��DI�vCO��q`q|��� �`
͂I��A.!�3���@�e���8��pC���Q��o � @�ME?Q�"p��J�g�T��P�T �Lp� ѝ � .��8�,�T.��� $DUMM�Y1�a$PS_6�@RF�@  � s�m��LA� YP9c��� �$GLB_Ta��Ũ�Г�C�&P�q��� X,��!�ST��SBR�� M21_V��8�$SV_ER�0O��p���CL����A�XPO��w�wpO�� �� D ��OB��sLO� I�6��\Ӧ�6���qSYS�6�ADR�qw��T�CH�� � ,xI`/�0W_NA�Ac��\uSR!?�l `��R p��僆�閂�塇�� ���㿉'��'��'� �9�S�.�9�w�ECX� �"��e��������|0�`qXSCRELj:��(�� ST~�)�}��D���`p�p_�pA9�� T,	����q� �P�B�q�A��Oʐ�IS�q���`pUE��� ��!����yS*��qRSM_�����UNEXCEP���{�S_�Ѵ0�3	73uCO�U?P�v 1��UE�����\�PROGM�pFLަq$CU	�POXb� P�I_�H�� � 8(A� _�HEB�� ��RY ?��d҂A�b�jүOUS�@ �� @��'�$/BUTT$Ryи!COLUM#��V�SERV�s�PASNE�p9����� 'GEU�q_ F� ��?)$HELPe%��/ETER)�'( �(2��(p�)p�)0�`�)8��)@�t IN� ��� NS �p�1�q�@  �vL%LN��� ��rw!_e"�$HB0�pTEX�sM0A1��^adRELVPDl��as0E5p3MV3?�,�5S3�tq2�шc��USRVIEWN9�� <���UН@�NFI�p�0F�OCU$��0PRI�[pmc�K��0TR�IP��m�UN����� ��B���WARN��� SRWTOL���	 5Q�V O��ORNVGR�AU:YDTnI���sVI����(���yPATH�2yCwACH9cLOG�G�ALIM���C6P���5gHOST���!�¥R_OB�OT��QIM�G ��S{РpU �B���H����0VCPU_A�VAIL���AEX�D!�PMT�G~R�G�{�N�``a�@�b�9J�2�a�Ev���$BACKLA�S�@Aq�Ab:�� � ��C7eV3@$�TOOL��$�A_wJMP� ��T� �$SS��Yt>`pVSHIFCP���P%�y��� j yRjhsPOSUR�s=W��RADI�1�d�_�ӡe��q�P����dLU��$O�UTPUT_BM�QmPIM����``�ܝ��cTIL�gSC	O�b�cC��d1B�f 1B�g1Bv1Bw1B"x�D��te~}R�W��t�Vy���B��D�JUUA8!d��WA�ITx�B�U%�pNEa��YBO�: �� �$x����SB!�T;PER1NECQ+�@?�'�� O���S1RY@@g��c<��$�B���M��7!���b\�@��Q�OP�JMA]S� _DO����T}�D@ m���0}�>�DELAY���JO� !���ԣ&��s��0���`��QO�\�Y_�A�\�v��c�Ah�$�? OaZA;BC��� �P����C�0
  �$�$C�P;P����ё{�ÐڐƐVI�RT�1ϟ�ABS�a�1 ��� < O`%�7�I�[�m�� ������ǯٯ���� !�3�E�W�i�{����� ��ÿտ�����/� A�S�e�wωϛϭϿ� ��������+�=�O� a�s߅ߗߩ߻����� ����'�9�J� ���AXLMT=PJ����  �\�IN8e�w�[�PRErP1P�j�����LARM�RECOV ��婀F ��q   dJ��!�3�E�S����v���������, �
"���V�NGXA ��	 =#��
+ �PPLIMCX?��Handl�ingTool �l 
V7.7�0P/53 ���
�0_SWq�
F�0�� 154�2��v�7DA�7~ ��
e��{:	lNone��m 2PO`��T�GX	�Z�P_�!V��Qu�6U�TO��;@k��Q0HGAPON�d��zQ1U
@D 1��� ����S�Q0�`Q 1�� � �����	�6/G%��\#֒�ܒ �`+$�H%�A*HTTHKYU/ג/*/</ N/�/�/�/2?�/? ? >?D?V?h?z?�?�?�? �?�?.O�?
OO:O@O ROdOvO�O�O�O�O�O *_�O__6_<_N_`_ r_�_�_�_�_�_&o�_ oo2o8oJo\ono�o �o�o�o�o"�o�o .4FXj|�� ������*�0� B�T�f�x��������� �����&�,�>�P� b�t������������ ��"�(�:�L�^�p� ���������ܯ� � �$�6�H�Z�l�~��� �����ؿ���� όZ,�TO BTDO_CLEAN�|4��NM  ����*�<�N���_DSPDRYRL���HI`��@�� ����������(�:��L�^�p����MA�X? ��Z������X�ā��6PLU�GG��ǮRPRUCs�B������ĝ��O�|�4SEGFzKX�j�u��� �ϼ�������<�o�LAP�߬�n#Xj |��������0uTOTA�L����uUSENU��� �ȋ����RG_STRI�NG 1r
��MkS2�
�_ITEM1�  n2��/ !/3/E/W/i/{/�/�/ �/�/�/�/�/??/?�A?I/O S�IGNAL��Tryout M�ode�Inp��0Simulat{ed�Out�<OVERR�п = 100�In cycl�5��Prog A�bor�3�}4S�tatus�	H�eartbeat��MH FauylGCAler$I T?BOTOfOxO�O�O�O8�O�O�O ��� ����O5_G_Y_k_}_ �_�_�_�_�_�_�_o�o1oCoUogoyo�OWORx���a%_�o�o �o�o!3EWi {�������8��/�PO�A U��k>�x��������� ҏ�����,�>�P� b�t���������ΟP�DEVX���l�� � 2�D�V�h�z������� ¯ԯ���
��.�@��R�d�v�PALT ]���ow�ſ׿��� ��1�C�U�g�yϋ� �ϯ���������	ߋ�GRI���Aѵ�� i�{ߍߟ߱������� ����/�A�S�e�w� ����/�iR]�� Y߿���1�C�U�g� y����������������	-?Q��PREG��� ��c�� ���/AS ew��������W=�$ARG_��`D ?	����8!� � 	$W6	+[L(]L'�W7m)�+ SBN_CON?FIG 8+�1��2�!CII_SAVE  W4��!�"+ TCEL�LSETUP �8*%  OME�_IOW=W<%M�OV_H� ??R�EP��R?%&UTOoBACK� �-�FRA:\�w Y?w� '�`�0w�2�#�?E n(w�?O2Op)O;OhO�4���nO �O�O�O�O�O�Ow�O _._@_R_d_v__�_ �_�_�_�_�_o�_*o <oNo`oro�oo�o�o��o�o�o�� � �1SYSUIF�.SV ��KCT�L.TMP DATE.D��\n�\�a=INI��w��%k3MESS�AG� �q�!@ �{ODE_D� �&�6�x�O���k3PAUS�U�!�8+ ((O;"U�g�Q���u� ����Ϗ��ߏ��)���M�;�q��0�:�TSK  @��?��n0UPDT�p�wd��
�XIS� U?NTE 2
8%�# � 	��'�R! �O�:�s�^�������p��˯��MET��2�Pܯ5�دY����SCRDCFG� 18%B! ��%�"N���Ŀ ֿ���ϛ?�?��T� f�xϊϜϮ����=� ����,�>�P߻���'#q1GR��ސ���_UP_NA07+s	q4��_ED�p�1��
 �%�-BCKEDT-`y�/:	�-����5P��r2��w
n"dOw����2V�.;|� ��r�	�J��
�y��ED3���g�����pC����/�ED4�� V�z�����R����ED5B�����p��ewED6� �S���/�	ED7�B�f��p�>/��ED8./�/2���w/�/Q/c/ED9�/�/??�/���?�?�/?CR ����?�?-�?(O�?��;����NO_DE�L�ߩ�GE_UN�USE�ߧ�LAL_OUT @��t��WD_ABO�RNp�N���@ITR�_RTN�w��LN'ONS4��v�q�E�CAM_PARA�M 1��
 �8
SONY �XC-56 234567890��� ��p @����?�H�( С�>Z=�F�]U�f^@UHR5SS=�vѕ_Χ_R57�_�UAffjZ@O0oBo>Ofo xoSo�o�o�o�o�o�o��o>P�zCE�_RIA_Iޘ*�PF|������=��q$SGP 1]@��~uߐ��#��{CI�D��F�PC�pC F�(�F�SPC8F�@F�H�F���CXF�`F�h�F�pF�x>��� +C�F�����F������ɏӆ=�jQPHE>�0ONFIG�O��G_PRI 1������}�H�Z�l��~���������KP�AUSPOS 1-[ ,E��� �,��P�:�L���p� �������ʯ���4:�ВO|���ȾR�NDET_V�2���C2r1KV��`�r��l���PV 7�ܿ�y
 y�￷q) �;��<�'π��;Y� k��Ϗϡϳ������ ��T��1�Cߜ�g�y� ���߯�����,���	� �t�?�Q�c���y�?GRP 2���r� i�y�IO q���Q�w >��F�X�j�|���F�}�TMR���'�
�E^�_MOR���|� �� 	  	,P>tb��D�s�����A?�큠��pK��R���PV���j�a�-�/A� tp����u��tb�w�i��hvPDBX� �\���
mc:cpmidbg�HO##:��q���p�U/> #  ��p�F­����/d*�·p+w/C/�/e)�D88~(g�/+?�-'?�f?s?)�u?�DE�F ��C)��b0buf.tx�t�?-�?� _MC��!�� �d,EC���"���VW�{Cz � B�q B��F�B�8�B��~�C� Cޢ��D3�u�zq Dz�l'D:�"Dr�BENNE�A7EV�ߓMF��pgF=C�F��e,G���Gp��G�/��y�jT	F�$��4Tm��p(T~�p�p%�G0�VT3P���Ag/  TRy�D�VP�a  EY�E� F*� F|�G�$ˀF[� G�R�k^Gl��G���G��&H���G֓�H���C��  >�33 ��AN�  n�q�@�B#5Y�Udu�A��t�=L��<#�
�4�1�o'�BRS�MOFST ظ>�rIT1<@DEg %�l" 
 av�q;�`  0o�*oNTEST�2#_oksR�r&\�#^FECPA�[偑�aHoBՁy�B�@x����S-�btT_�0P�ROG �fr%��?��vINUSE�R�铄vKEY_�TBL  7���Z@ �	
��� !"#$%�&'()*+,-�./��:;<=>�?@ABC�0GH�IJKLMNOP�QRSTUVWX�YZ[\]^_`�abcdefgh�ijklmnop�qrstuvwx�yz{|}~��������������������������������������������������������������������������������͓���������������������������������耇����������������������ё�pLCK��|��s�pSTAT��s_AUTO_�DO  ��F�INDT_ENB;�bw�R�aY�K�T2����uSTO��~�R�T{RL�pLETE��� ޚ_SCRE�EN FJ�kcsc 	R�U�ϐMMENU 1�'FI  < �|�l��K�u����� ����毽�ϯ��� R�)�;�a���q���п �����ݿ��N�%� 7τ�[�mϺϑϣ��� �����8��!�n�E� W�}߶ߍߟ������� "����1�j�A�S�� w����������� �T�+�=���a�s��� ����������> 'M�]o��� ���:#p�G+�_MANUAyLӟ��DBCOu��RIG��$�DBN_UMLIM��,A�u
�PXWOR/K 1(FK�o/�-/<oN/`/r+�TB_� )}��Y@|$�_AWAY�%�AG�Pr=�`�&�_AL�=��"�Y�Ґ��p�_�0 1}*�k , 

.�:/�d2?o?�6� M�t�IZ`�,@`�3OoNTIM��t���6�)
�u3M?OTNEND�4�RECORD 1�0FKUB)O�1�O�?A-O�k�"kO}O�O �O8H�O�O?O�OcO_ *_<_�O�Or_�O�__ �_�_�_�_�_o�_8o �_\ono�o�oo�o%o �oIo�o"4�oX �o|�o����E �i��B�T�f�x� ������/����� ���>�)�7�t��0p. u�����-��۟͟� ����N�`�ϟ��o�� ��)�;������8� ��\�˯ݯ����;�Q� ڿI���m��4�F�X���"TOLERE�NC�$B�	2� L��ͰCS_CF�G 1 ;x7d�MC:\��L%04d.CSVYϲ0c��x3A ��CH�z0_?x>��Gߠ}<��RC_O_UT 2�+-0�z?��SGN 3��%�2��#��12-AUG-25 17:24��O27-MA=Y��4:38�]� Z�t������x>�з�pa�m��PJP���k�VERSION� ��V2�.0.11~;EF�LOGIC 14^�+ 	TP���P��p�PROG�_ENB�/B��U�LS�7 �&p�_?WRSTJN�0���2�$EMO_OPT_SL ?	�%�]�
 	R5�75x3?�74D�6E�7E�50i�d�o��2E�T��j�"�TO�  .����k�V�_�0EX�d�5� PATH A��A\��M_~;�ICT�!F� 5� 7�$`�e�g��}STBF_TTS�8��E�3t`���MAU�\��2MSW��6 9���}<tТ�7�*! ��]lR�v������DSBL_/FAULy�8�/�3>!GPMSK��2�TDIAG 9؍��`����12345678#90x'S�lP���/ �/�/�/??%?7?I? [?m??�?�?�?�?�?�L#@PV/ � �"�/�� 2OXOjO |O�O�O�O�O�O�O�O __0_B_T_f_8Lx�gUMP$�I� .��QTR>;#�_�PP�ME��_Y_TE{MP��È�3��84���TUNI	�w��YN_BRK �:��x�EMGDI�_STA	���GeN�C2_SCR ;7k�/�o�o�o�o �6�o�o 2r�ncUa1<yo+O|��в�lbTt=7k�Q������o>�P� b�t���������Ώ�� ���(�:�L�^�p� ������ Oǟٟ�0� ,���+�=�O�a�s� ��������ͯ߯�� �'�9�K�]�o����� ����ɿ�����#� 5�G�Y�k�}Ϗϡϳ� ����������1�C� U�g�yߋߝ�׿���� ����	��-�?�Q�c� u����������� ��)�;�M�_�q��� �ߧ��������� %7I[m�� �����!3 EW��{���� ���////A/S/ e/w/�/�/�/�/�/�/ �/??+?=?wa?s? �?�?�?�?�?�?�?O O'O9OKO]OoO�O�O �O�O�O�O�O�O_K? 5_G_Y_k_}_�_�_�_ �_�_�_�_oo1oCo�Uogoyo�o�o�o�wE�TMODE 1>v'Ufq ����oGwRROR�_PROG %��j%���HwTA�BLE  �k�1_����jRRSEV_NUM �b  ��a��pq_AUTO_?ENB  ��c�Zt_NO�q ?��k�a�r  *U�6��6��6��6���p+5�O�a�s��H�IS�sXq�`�_A�LM 1@�k e���6�6p+t������&�8�J�x�_\�r�  �k4���b���`TCP_V_ER !�j!6�Z�$EXTLOGo_REQ������SIZ�ܔTOoL  XqDz����=#�
ޒ_BWDo�%��vQ���w_DI?� A'U���dXq r[�S�TEPg�y��`��O/P_DO��$�p�FDR_CFG {B���?Zp�A   >�  �@��أEATUROE C'UQ��a�Handl�ingTool �7� 5\rb�English �Dictiona�ry=�605.AA VisS� Master0��>�0iB/a�nalog I/O7��>�PRINa�ut�o Softwa�re Update  B/16���matic Ba�ckup;�duc�t��ground Edits��  D pr�Camera��Fމ�1
P�el�l��ʱ7in�o�mmj�sh�8�87\hi%�co��=��ct\h%ǡ�pa�ne6� R J8�%�tyle se�lect>�\im��on߱j�oniwtor<�h73x��ntr5�Reli�ab��<�0y�Diagnos��䂱:�
����ual� Check S�afety UI�F z�1E�han�ced Rob �Serv��q o�Ͱ�User F�r�>�A�E�xt�. DIO ��f�i�� #�=�en]d�Err��L�\�6`�[�r��C� �@�:�IF O�FCTN Men�u��v��>�g H~��FTP Inp��fac��?�6\a�Gذpl�k �Exc	�g5�Y�High-SpeзSkiƳ  ��!�)���G�mmuni�c��ons>� M=-��Hour��p����R Hx�����cWonn��2=�(��Incr��str�ΰi�<�
TE�KAREL C�md. L��ua���pV�s�Run-�Ti4�EnvU� �"Tq�z�m�+��sn��S/Wɲ
 �License���'� L��ogBo�ok(Syo�m)���oadMA�CROs,��/O�ffse��art� ��HG�RÊ�\a�p`�MechStop Prot���d� \h64��ie�Shif��9�鳇MixЂ�����C�VL��ode S�witch��c.Mp �Mo����.�� 72l_����g�'�l�!��ultGi-T�����!W��Pos��Regi�o���d#�Pr�t� Funb��II9)��NumЊ�>d� .com12П Adju�:�4�1\LZ� J85<P�ktatu<�wmm7$�RDM��otN�scoveW� 44Wѧ�����uest 7n�u`��oGЍ�<�.�fd��SNPX 9b�⊸50S�[��LibrV�'"L�o,� S��P�a찠�Ets i�n VCCMa0�ѣ� ����Z£��/I����TMILSIB��7eP���AccٰᵹTPsTX"��0iCe'eln��r�e�4��8�O9�Unexcept�omotn��  UЀ) -�7�N�f�� Q
��a& t�Ha&SP CSXC9�`����%[�3� pI �We�'�^ \��$vr��	�men�S  N�iP^�ax �
7Grid�play ����6�pŴ��0,�LR�l���2���%K�Ascii��l��7��v��st1Pat��6��OR�yc���� ori��� M���7ata�qug�c� ���[�,�0-��ЛRLEam��$5~��HMI De��(��� 7���C�߇�	 ��assw�ord?�L% � p����7�"A Y�ELLOW BO��4ArcV viYs����IF�5t���OpA�;�s���spk 2۰a��po�1 ����T1����2� �HT��@�xy��"V'���llig�� !Q@@�� !0�JPN ARC?PSU PR\<��9��OL?@S;up�Bfil�0Z��2C!uQ^�l�cro��mS�L4 ES�T�SS?@ee�tKex^� J �Qo��=t��ssag��@��mP�P��]�!	6=2_�Virt����9�z�1stdpn�6���SHAD�@M�OVE TF�MO�S O��45�get_var ?fails ��o`�%�AE۰�� Ho�ld Bus$$C�VIS UPDA�TE IRTOR�CHMA@$�iWE�LDT�S st��Q�a: R741�-�ou�`b��62��!BACKGRO�UND EDIT} Sb 26.f� �EPTCD CA�N CRASH �FRVR A/R�@�cCra.�s �2-D��r��$F�NO NOT R��PORED �p �.pJUPO>0 QU�ICK�`OP FwLEN�Loc����bTIMQV8�F�PLN: wW��p�lT�FMD DE�VICE ASS�ERT WIT g823`�s�ANTq�ACCESS Mv��JoQui��p<�|r��x�USBU�-�t & rem�ov��,SMB �NUL	@lqER �FIXG��HIN�]aOL�pMO O�PT 23g `O�ST?@wDU h��p�dAdd�adl.е@io � AMp�P�pWORD.$�apO�IN;�50��aP:fix C�PMO-046 �issue 16���J`qO-P1�30��TES�dS�ET VARIABLES^`����c�3D m��vie�w d(M�W�e�a��8 b.�of �FD ��л�Px� OS-144 ���h s c
�p�t�s ��lco �� �hWAp���3 CNT0 �T iLB�T�I9m��Z�ca mq� �POT:When���ews�STY �M120a�t��p�t|ado GET�_�� �,VMGSR qAWpA�@C�a� Pq@�C@�ͱ�� �C�@� ELECT�?�L<�ING I'MPRPQx�RY�\`�s�PROGRAM�OP�@� IPE:S�TARTU�AI�N-l�  ga�S�CII�`��OF �LO��PTTB:� N �MLK4me�0��:��moW�a�ll�pR�L�8l`Tor��AH���yS1�QP�th�pn�P ch -р� yTU@�Rtou��5�iR�Cal��Sig�n� P��xUThr?esh123$W��Hj� : MSG�_P4�\@er  �ap�G�A�ze�ro5 ���@ 6t�c�d:��U@��2Dv� rc�OME�p��ON�`f� 0;ASREG:wV^�őHt�˳KANJIصn�o̐0Аc�@��n� d�1�QTEQ�IN�ISITALIZgATIpD�Awe��� =�dr\��D�c���minim9 reAc0ˡ�c@���mU�?ro  iC�dϰ=�i��({���vd=w�� 0iB�Ѓ����w u-�mse$SY�`M-��q0�#%�bW�lu��dӓRe�eÂ1T���m� t06�0War�nő@�בBox �fo�PseqPVEORWRI�`��S��ڿ�F��up�de/-relc0d"��������őbetwe���IND *��igE snap���usősp��FT�PDT�DO�TqH�ANDL   �Q�d���D4�n� � D=����ope�rabil�0  sH5�[�: H52�0l��ܲ51�!����mp�qs  Jk52��O�pFA�P|_�^aV7. )U���`GTH�pi�s�ݐ�0��mq���ne-RemarkE��� RM- tp�qtQfPATH {SA\`LOOS���[F�0fig - GLA eli�Є����p'�ڤd �!E�ther��� T�rac�� H55��W@r7O� 2
PE���>�80In�P l\0Q:���Ɛd|�y��it ��P�p��Pay�1[�2]��
�Xe1:� g*�s��dow2Dt[ �@IS ����EMCHK EX�CE|�1H�MF I+���qh��PnHPZ�P�qB��Ĵ��DXr�8�0 ��c?�α�e A��E�Fa}l1�alarm�� V��IRx`[��av�1�r��aopX�� ck��6pr � "y��@������Stud>��`b� fp��: U�0B�UG?��2��DUpP�ET<���� �S�E�XPANSI��D3IG+�KPO ��dCCRG EN��CEMENT �p�HM��K ���pH GUNCHG�`�EXTEpP�c�
�aS� 0q�����ORYLEAK?���4��pLC WR/DN R1�O'�
N��SPEn���G[�V *�|!MU�=�7.�SGRIHA�@��0\t��MC E3TH� ��SUh��p� 8Y��PENS��`N�P8�[`0a��B�ROW�pR�RMV ADD ��rA��DC��pT3 A�LAcP 2��-�V�GN EARLY �b&�����wr�!�LAY{�8� SP�D��[PHM#S "�T1�0TOUCHi��Ї�F��JaY�y�|5 _ERRORF �DE SA/<@W{RO5�CURS� i�I�N np| @�[!-158�G���ORSR �`TqU��(�7@�6T�"F7�"@�s�%1�%�u@!B� SY RUNN4��9�p@�BRKCMTARO�dP �@�`AX�`��PƐx��@��ISSU/3��C$pTSI�1K�WCIPSAFE�TY C(ECK|�59=#qA4�w0����=�� \!TWD��R41ǱC!INV�-�D ZOP��R2�4;%z21DUAL�6��ӁC!S�FT�E�� b���!0NDEgX F� �% X���%UF�BP��h21�!�4RVO117+ A	pTg� �PT��@�FAL"TP2[47�Rt\SQP[An�HIG� CC���SNPXF MM �!4�@��t��V>�\���2`�DETEC� `p@�� "RU�K2�PuOS5��Y�6@L��G�� �vWT� �� 9691�U� ROPP�P B~FITP4MS��qgkϑ@�RCO�PYG6IA_�[ �T�@4K�`�6IA"�GC�U� i� �`A� SIZE 67)4�`O�7��-\0��!F_RO��D�CP� PA��pANUC�؀S�IL�.pc�` �`RE�s��pl�e��  gtpa� �`
�a�����\r�b���utal�a}p�`sn	p '�1{p vKt21up�|Kpcir�b� JqslDqhtp1x1!spngi���Cxkey�})qgvp1m0zp�|usu!u]g-�.vr*���� b��s�]��0�$q��~�!! j921p���pl.Coll�	�Skip��y�R���J��*�3�� ��il�q�� (��, x�A �Ar v��.��]~���>w21\a=t*`7 "KF�Q��,����\tptc��"TCX�m1�}e�>pkmain�;�setskck0| ate�m�s�F��郣�Y7���KA��U2 {Sp��FCTN��H�0ЀpJ��ڌgՀ=7��AREL�������7A�����)�(f�)q*`8I�8O���Q�h�D�9I�9Q��pz�k���rp"K�RCF��s�ڢc�tme "CTMqEO�Z�أrcf���p|�(�!���g�pcfcstmT���,�cdt����+�s��r�pb��ٖp󖦅73�P��p=�� ���c J�$��q(K<� � N�p��m�p'� ]�p����?�b÷�p r�c���U�寢rp�� �9���,���Y� ��q v�_���p��̑��̲��q[�й���52�Zd�C� uh S�et
  ���� ��J	�p	   r\�tq_zmove|o׹�finde�ornt�`�Ѽ{4��p�L�p\fnd�rٙ! 4�r�t�cpmate��T���M����0R63?8 R517˂)����(��aDqP�	�t�(q��m�%�����B�99��8�pp�,�i����p�PM��)�etg�uid "GUI0@�y�V���spe�)q>.�tm_mo������refB���a��8)�)q��log�P��prmpA����va�(V�������������	��mas�k��Gq��sk �Exchangex����2H541%�93*0%c�96H%0&9%B5)Dp?2��1��u�N��v�m�x� ��0�I�0k��t� " �1£�}��H���|�Y�dsuch��P�sDi�yIm�"�v҂8@�&�8�87 (G!]�isplaT%��RƠ]��9%�x9 p�"*`2RI�2O��+t9 c�D�@x�� ar� 9&���(1sca2��*m��scrL�BsX8trld��S=��9(��p�8A$ayl.��`n�firm2#b'78 ڊ��A�  K��@T!��{8B�3I�3�/�]Ei�plcf "�PL�?�Dpfca0�8\�A���̧D�Bov�?Yin1im�~V.vp"&�aA�r6�A��Sh�ape Gene7rat��IIDQ��c74ڈ�r�R (�] p�(�p�a�^|�;���K��^�enuu\�hD`n�HMN:A�;cgil\D`<`sug?cia�nue�Bshf i���fhi �Ofd�!��tm�?��fh�a1vY�$|2�o�k�aq3<�iodsm�;jenR��7mensub~~}�fh� �w�$yseQ��w2�crc�MSfhst0 H�kc�Q6d��>lbdetbo�k� gk%E^fg8�
p����	akadspweb ��Vo�x����S�8��G�:b201��Y"|�3�����4���9d�5��"'e|�il��@����[,���HA���� (CalbP�,q�_aca=P�_	W@�4�6;�6��؛�ţU�mt�LM�T�ͽ�et@��A�Lj�-�몶��7ţmac��K8ån�sv�3����� Q����c_��@i�~Y��joi�@�ٟ��F Y��_trc@:]�o����c�������0@���4��}UCenter aF5��1_�20\0{��ɚ&)¨*4�(�/p�5�7;�7�q/�� "F���.� ���;%�4��������.��qp���W�a{��g   u�xra�paxr'mrf�oG�x��"&�K�/'turbsp�ed�T����W015�P2�����s)��(��ya�_�F�⦯8K8��P�k97Т��|�$�1.�8K�788���'�tsp���1�?"���glfmԏy�st��&�R0�O�*�vr����� vQ���@a����Y�| pshi�m��P�Pim (~xTool)T�6������ ���Ale��]q��	�5 �B�fx@a "T�PSH�s'pe��FLEX���' 1�5 b�R�R�r�%B� l�rE^P5 2�Aѐp����p7adqG�DQ��5 �]�8K{ �A4@DQ �_��7!	��1s7�!/��95��+�1qvl "DQVL�	d�$�dq�I�I�&c3c�  H55�2_�-121 !d?AAVMS-2�0QpaE0TUP� s�J5495o�i0616?0� VCAM @R�CLIO�#gR6m0� dq�0�MSC{c�2P�#STYL r9 �vu128@+��0NsRE/#�0SCHS�DCSU r�mal�0ORSR� c�u104��EIOC 3�Q��0542 ��@SET Easy�0�J5y0Uk`(i07�y0��MASK� ��27#�0HO'CO )�5B3�Ci2�2W�fik5B0 �8֠#u1U0p553�9_F�A"NORM�LCHKK5O�PLGQfii10q3�0�M@HCR�RM@C�0aAf�B6���i154wEMDSWBuQi@���137��B0�Av�@7@PL+��C7 ��5B53�N5B7  <A�B5�S�PRST 7�7a�FRDM?  J989�0�1���-0930�R�PS�NBA uhQ�0H�LBGESM�PTDS'PVC#si12V0�-0TCP��T�MIL��PPAC� k987�QPT9X{��PELN�c�B�97�UECK� L�88-`FRM� �� �1OsR 8�0IPL+U�CSXC e\s=w�0CVVF�QKTP�Ad�@��6O�rob�0Gy`��I�Г5IPGSns-08%`���Pz��7eR663�p�se0Q523 "�rkey%R1K5Rw696{g51 �a�.A53�U�01 :~`sh31 a��4A�6%`�AA75 t�� �0�`6cal�`CTOP[�A�0>pc80 sler�@OPRXY�57p0v885 rec;QSOL�0L4S}� q}e�0LCM h���lPETSS��%R6x��`�PCPE ���PVRC�t�bN�L�eU002 uĉ3�p6� <p�r7 B�at�q�@$��1�ej�4�m�5 > �W\0U02"@se� CI�3sUK�4 3822rK�5 p��q�P(Wai��`R��o<�3v@��y�VU�046Po
��3 d�"��435��6 .�(�q10�A1ق4�Eۀ�5 ac��ق7 o"MCR`�61oe��4�AmH�65 S96J�	�6��PT��68Ǉ�qpa�7	3SuG�77�qipM�&̂83�5k�4�"<�"�pw��pk�8�Uk��9����q90 w��s��1�9"@��9�5 f�u97�5Uq15P����101w��vFU1M���H�1�qP���7 ���86OP b�PU1�@=!%BA�1OR$�1AQw��6�P��5 16 (L��`o"�NPx�푡Pt\bu<�1�`�z��s���`��!@bbf��m0d�Ǡ�fU1U0boxi\�`�1�68,��1P��58��596`69��60ק�����p'�6 B7BOX �67�u'����psche�7�1[�72g�6 setu����\��p��ޝ�offsH�93�K5ð�b?�2)�btcas�@۰��21��219�Pld��2D�`��2q����2!@'xcdg1�8o5��9 ���2U0liD�E�23�Ep@�55P$ ��� =�<�5�p�4k�3 or^Rk��psro'qk�6 y���i�7 �i�9[�R�$��A����2 P �Eoq��6 very,��9 ��i���ʃ5q� ���8��5��P ��`��5��9W71"��3��5��re��!@ecj�a O�
@��i��`��	pK�q�ƀp�p�8������6 ���7 6�29 @@U5�pa�nagH�5����57��5��*`�a���7>�57��Մ58�2 4�5y�ĕ5���o�i���"XRM�@?�2 C  ��=�3 	�K�	=�4��99#�6 �@�y��@y�u@d�]6AP\acׂ6��Pe�y��0ĕ6�Pvt�z��6��"ACS��7{�6E�_0�qc��0�q�\�9�sv~�`ANRS e�r+� vs!�h���~Norchma��3� � =�Ma!��!�� 39 J59�!�598 J68�1 !�7e�`J6�Q�W%!��c�!�L�te,t�s&!��P�#��lA��� �$IF!��AARCRt�1 �H��a�o39�:�\9�cp���P��s8���FA!�H597v��92!�LSE�#p]�[!���tmk]�64`60�A� ��F��t�1%�!�&!���or!�S961 !� �!�kZ�x/0 i�!�9�?���f_ �!]�!�� !��4��)i���(��tm��]>�R�h�����A� "TMA�`�&��y��in�_!��A��Mp��!��&����et�d�2���&!����moveto��%���?�9�mmonitrD��&!� �T�onst,"��a� D"YDP��^Q�! paraHI����ame]�Cont�rol8�W�@!�4�3`�0@^�25 �R0�588�P0��`��t�]�� (P�P�eter�"!�, ������R,$�"L�Q mB�;33�� \ �E/93�ap���e�2�� m2�oladjk.f]�T=p F�2�AdjustA�1 `��18BZ81&A�J (�2��e �3�$2��e02j�2\P�E5`*C,�;adFADA�V
�� .@t �4��m10s>OPGj��O+B��p�	!	��1�#8��`��^PI�!�aeP�1aBi�3��N56�3 H]�(D�r,�ol 4Y,4Q%r���ᩢbLaq�r� �5 � !�.<r�E}C!�������vC3Sd`!�f�i��PFI`NyXsltpal�_�Z�tpts�TSR!N�[�{S,�pf`
 �sw�\�� ��J	!�	 �  ��J-RSe�rvo Gor@�������u'j���bT��fD[����j6�70g "SV�G/`Q�eQ%�aA2py "CO00qX��, 0��o�fsgn "FSG Q"17P.�`sf��XaPSW�
fB�A�e	!sgatu6p!�e���asgtp!TGPDR0o��bs�19�79o3�(sPp��t,��`GATb�Osp!�[sr*�bsgk95*��WYq?�ftdL�ߐ����<��rtdfl\!�<Jځsmchh/b�tdmen�2I%�m�kpd�1���xhk�wmvb�󈄐�ku2�f�mkl�w�0���fscli�ni/)u,�ldv	r�"�v�1�X�9��J�,Q����`�aaut�p�7A�S���1re��sub�'P!�Nt9 �aZq����b4Au��Muh�ĥ�hk_�kvP�Y  >�Yq1�P�H1�|ف�tol.p1� i 1�7�H 1�G��`1��sev��1�g� u 1�w�K 1����`1�kksk�Y1����, 1����1�Ƿtch1�q*�$�1��p 1���E ���uk݀�� $�v�1�'�Yp1�7�H 81�G��cl.�d�0!�t�1�F�\j1�J��r�a���1�v�VL�!�Ĺ1�gtsgvaٴ1��q���1�Ƹsg1�ex�Y1�2�0����pr1�7�gcre1��
I1�f&�571�6�du1��bf4p�A������B�0�E�%��a.f1��B����� �cSch�e��T���Ho�44B� 8P1��%��S!���d+�1� 2  ��H� 1�	�Ktb\q��tp��0b0�l� ��1��D+�trackin��0�����P����enc �01�����q�i�K!�1�������alts�t� ��E�б�vr ��1�e��P��ם0�Ѹ�41�sba�CV7ers1�ll�Bk���!S� �(Q�"(V.��Bel=UI��,6}�baaUH01�u��ssT`E`�
d��$��b0k�j05��sb��9 I�����9��F� ���B��en���C��(QDevices��:�K�����|�41�86 (O�P,�q�es 6)�@P��aU$A�o�\p3k!�j1�p
bx��@�Zaopn��`����|�1�pc��䌔��o`��glfm_���V���&���V�sc��a����~�vropio�@ q��E$1��A,�1�)p@�����818�C�NEM��mp��Jx� ���! (NE�ump��zǴ 1�XF��1nmn�6��SeD1�42m��T`M�PTP�RA� 61emocol���33�mpΐ���"�j�536�A1�uch�$�ns�0p1��J5Pp���$S�3T�4�1�ngP% !60p1%	P�36�d1THTK�1Dq��0�\etth��TH�S�sJ11*�01�hp�gio "PGI�O"PEp�vCth7wkf?FMc�ƷMHC5�48�5�2�V1�xAmP��q5i7c�� �F51/��F
Ttsn��SNSx�����A1�8V�A8q?SA[Quif��Q���*�xAp@�t/uD�A�M0�6X5 Ѥ��B ^P�ٙ(�2�	��Ѹ� �dQ!�`��1RJ؀E�xN�y�1� ��J��1�ipc���ݥ` "ctsk�e1*�`�R2k' ��!��a��n!�acc�0op�4�pC
p���R630��aX�)p��tt�!Q) "q�u\� �:DJ3��r��pawachZ@ACH���dOfw`�4>0K94�D3AO �u3k94����p���q���chflo1�ST-�v �/Suq�h��fp�A9�st������w�l�)�sA�?chcal2L�^�6�s��@�F�_�%I��[�vr	r�jv1�!� pai�aQ�RA~��Waterb@�,����56��L@����5=0(t���}�rnet�!QTy�$j�5B���xv��ؒj�aICS8k3o`�\p4�p�t �s���&�1��p�w1*��k�ta�`��k��cc����D���cg#en^����cf���C�Ԧsp�E�Кpa!w����ؒi�c� ��O"D���ѱ��q�Fgԁ!�w��A��ow��!�R50�@�3��,��ư (0�F���/ *���5C�q4��$q� �r�x!�]P��Mp1�Z�55dA)�ð�ѥ�*/|�af؀b����U�a�i���(���af��|�ep�0��ca߯����Qh��Ҙu���2! ��L�ine/Rail3 T�䷽69ɿ�� (�����FWq�i��0g5OGJ��p8B�r8E7��\�9�r`�0E	�%��q53R=3=� ��f�aldebu���RSkr���q3R3RzA� ��pgdb DBG2X���!
�H��ۀ�� ���2Q��% k�Ѹ����`���MH_bper O�ption�c�78���	P� ��`��0���Z'hg�`9Z�m��ht_3F�q�mЂ3k�At��qd8iᏣa�9����et�w��1 Fb�pl�u� -�.Handl��O�q��&V!�-G�P90�P7�A�9�Q(Ma��A�� ��0Uy�ܟ.�fF`138��F�!� �hH�qE?���x u!? ��O� G��"fhnd "FGHND�!T�&g���wמ#�Ic��lio��#Ce0�/O�+CLIO�A1�񑑜 45�A9�C�1�4�R S�[R�AR�!J�JO�ELSaE��1���"(CAI/OG�B%H�$��O \c��G1��Q��55h��e0��tcm�ACMIpa4�d69t�a�0L01�1���a�2iomenu(?�qAf3l7pc 1���8��� F�xe2�d1te1+��9dt��|��7eFFd���bW`In�t 1l Pump� Cont� 䐑��a`1��4 (��A_"�Hl,����E��!�ha�quy���apa�y���5�q�r�q�?:Sa�``1PCD���n���e�`cnd(j��Rq�p��a[O�Q@ѣ�P�Q_���Pa$��� ��2k�� ��a��Srt���?�Q�Qd��b!o \  ������	   ���#��� �&��$��J517 (Pr�ogra�jus�t�����`�� j$rG0�0��Ds�1�j "PADJ����Frprgad)joAup�ppE�A/ �v���3�v`�f�Dp�1���j539`�-� KAREL Rwun- �Env����! J��#�13t���`R0�J97�!�"6�!�c�!�a�e��2�"�����F�(<2+�ime (6�U1qe����.j�p1klut��"U�TIL@#�\ewtqm_"MGR/ڄ H 1���11Cp(�kcmn���Q��J�\��sߖ�qq����ex�<M&�q�tr$�f�������;tp�psts�����a Statusr�+P�ѩ"H51  e�"v����g�Җ�зPR70(�17�p ��W���&�a!戀;%�Q!sHs2��y%��  ST�D RSC�LANGc5�أ5�?prscrn5��5�֣Y�.v5�i�5��+�5�dsblf�l5� Disab�5�lts�5���C 5��#5��ӡ�25���3le5���ar5�V5��ds5��5�U3�l133Ą�5���5���t\��"DF�LT5��=�w@sbAf5�����M�du��.a�i򹵝�j5530.��q P5��5�J��_Ÿ�5�0 /(Adj��nq5� 	S5��Y���5�zq���5�34��ݵM�E�d�q��Vs��Jb!�*�sh5�AP�5�J#��\a���Ra���+�@�SY�W�M��q�� �C`���4�'�p�ti�P
ĹR5�7�|��5�)(&���sk�,��R�RBT"�O�PTN ��� ���b��K923a"��d���0ol��gP1 ���������rcm\p��57���DPN����K�ccf[�J�I� �K�@,�K���J�h�J�o,� I��QI��I�l��I�s�I��Ӟ���I�n�cy.0�UPDTG�����o����� 3����I"������io9v 2byn���� l������Q���
����acc������2��p� 2��ɒ�� L�R����R������.�a������ ��Q�!�+-���� �������2���� �������� v����ex����	GcchW�F4	m�aq! �H�w!uTo��sq�!��汮��Ry&P �n���u-1�82�iag�&Rq �!�����5��q
�p�92�DP��) � 6SQE>���pi�t�G��
�pg`%p?�4mon�?z?�?��vr���?Dgse� /��f�aE4!  7�e�A�������y�F3�b�%R823�%lA�c��E4	R�.���5��Osl�k9�Ur��*FP2�6E48ÚsT&ed�g%�O� GVTD3G"%*sl3F��_sl��_�Z|`s��_�[�1�_�[fil O�\<I�-�6�X8e ��4�U&zKJ5ٲ�F3m�%5  �>E4	�K	�O/@����?��tstn��ƕ)pD�)pite ptoo)pƖMq���p)pErulsu0)p�v)p^ttl)pjtC2.)p�v)p�uiMqtupdcyc���|vr�P��x�1������N1���qt eq��)p�r)p�)e��3���o��P"�7�@q�4���?cpy�r\�dqil5œ`)ph��r��l6Ŕ )p�eq��pq7ŕ)p�����Dsw$�,>yx�f<�ǖ�]u�Frl�k2dq�*�conxC ��wcnvu����bagtch���palctr����slpğ�iOnit0"�4�mnp h�z��q����fя�ebT�iu��cy�R���Dsv<��𿯭�)b��s<�d����h%�ߍis�axis0�z�b�=A��Crmled\��w�p�s<Cz���u304�Կ�5���502$�.�3@��� �s��|TC��olutlF!�aam T�B�ox{�I�w�59m8�90�`73C�0�AӦ��� (�`)�� Q!��m�r�"0�g ES�"��sw�À`�Y��#F�����@0}�2�\Rc�Yxl� �|���q"TLBX��x�����olbx��tԩ�\t�ѷ��;� L�x��-!��-� Com�0��or� Cha���Т�F�h!e�OCM R6�14���B���g ��(��on�����?nge, P����BT��}v��*��B	��qr<�{xF�pak9=6�� 61R_PXZ���cr750�7� lV�h�22h�22~����Ѓ ���J	�	   �all<�mreg�!"J��?r�W�'�m <�����I�(q�R�m�����>s��5�=A}aF��'�.f��p¬q�aA,�l�qR  Tu�r����Eu�93 /J989h�9 �m�d�"�`�'�Q � ��+�i�4�E�N�|��p��P��X��Er���"MLEDB1� |����mk9530����8՝����YCS8SJ�\�ddqS���3re*��ip����&��igr�tM��@������>ydk� /*s�$/*S�<�H��  �D�� |9	�!�!1 C!   E�v�  ��# 	�!��"@�؞H�"  ?���E �8�� �P�<�*�gelpq�yx�"���'99 CP� ���$FE�AT_INDEX�  �# ��   50�ILECOMP �D���b1�P0�#U3SETUP2 Eb5�l2�  N� �1U3_AP2B�CK 1Fb9 � �)�"�?�? # %�?�?� e0�? )Oo5�?UO�?yOO�O �O>O�ObO�O	_�O-_ �OQ_c_�O�__�_�_ L_�_p_o�_o;o�_ _o�_�o�o$o�oHo�o �o~o�o7I�om �o� ��V�z �!��E��i�{�
� ��.�ÏՏd������ ��*�S��w������ <�џ`������+��� O�a�🅯���8��� ߯n����'�9�ȯ]� 쯁���"���F�ۿ� |�Ϡ�5�ĿB�k��� ��ϳ���T���x�� ߮�C���g�y�ߝ߀,���P�����q9�0P�? 2�0*.cVR��H��*K��q��w���2�PC������FR6:D���������T@0 @�R���=�|�C0�����*.F5�����	���� ��$��STM DMX����E���iPe�ndant Pa'nel���Hz��j��-��GIF7alM
���JPG��l����5/��
ARGNAME.DT?/���o \S//����$�/@/	PANE3L1�/�/%o �/?���/2?r?7 `??/?�?�*3�?�?@7�?�?�?HO�*4O�zO7hO%O7O�OK%T�PEINS.XML�Oo/:\�O�O�A�Custom T?oolbar(_���PASSWOR�D�O��FRS:�\k_*_ %Pa�ssword Config�_���_ �_�_+o��Oo�_so�o o�o8o�o�ono�o '�o�o]�o�z �F�j���5� �Y�k�������B� T��x�����C�ҏ g�������,���P�� �������?�Ο��u� ���(���ϯ^�󯂯 �)���M�ܯq���� ��6�˿Z�l�ϐ�%� ���[���ϣϵ� D���h���ߞ�3��� W����ύ�߱�@ߪ� ��v���/�A���e� �߉��*��N���r� �����=���6�s�� ��&�����\����� '��K��o��� 4�X���#� GY�}��B �f���1/�U/ �N/�//�/>/�/�/ t/	?�/-???�/c?�/ �??(?�?L?�?p?�? O�?;O�?_OqO O�O $O�O�OZO�O~O_�O �OI_�Om_�Of_�_2_ �_V_�_�_�_!o�_Eo Wo�_{o
o�o.o@o�o do�o�o�o/�oS�o w��<���p��$FILE_D�GBCK 1F����p��� ( �)
�SUMMARY.�DG��|MD:��[��pDia�g Summar�y\�iz
CONSLOGQ�4�F���ߏ�n�Consol�e log��h{�G�MEMCHEC�KՏ��J�c��M�emory Da�tad�lw� {)}O�HADOWY��>�P��t�Sha�dow Chan�ges��s-�?�)	FTPҏ?��ΟC�n���mme?nt TBDl�lw�@=4)ETHERNETa��~"�����n�Ethe�rnet ��fi�guration��spV�DCSVR�F`�F�X�q�t�%�6� verif�y allt��s1�p�1�DIFF�i�O�a���u�%��diff����"��6�1�Կ�{� ����ϭ�	9�CHGDE�W�i���u�!�&ߵ�9�2�����σ� �ϪߵσGDM�_�q��u�8�.�9�FY3�����ߋ� �߲�߃GDU�g�y��u���6���UPDA�TES.U�;��{�FRS:\S����o�Updates� List����P�SRBWLD.C	M���|�������PS_ROBOWEL��g\n�� ���W�{� 	F�j�{�/ �S���/�B/ T/�x//�/+/�/�/ a/�/�/?,?�/P?�/ t?�??�?9?�?�?o? O�?(O�?!O^O�?�O O�O�OGO�OkO __ �O6_�OZ_l_�O�__ �_C_�_�_y_o�_o Do�_ho�_�o�o-o�o Qo�o�o�o�o@�o 9v�)��_ ���*��N��r� �����7�̏[�ŏ� ��&���7�\�돀�� ����E�ڟi������ 4�ßX��Q������ A�ï�w����0�B� ѯf�������+���O� �s�ݿϩ�>�ͿO��t�Ϙϧ��$FI�LE_�PR�������������MDON�LY 1F�Ņ� 
 �5��Y� 0�}�=�f�/ϊ�߮� ��O���s����>� ��b�t���'��K� ��������:�L��� p������5���Y���  ��$��H��U~ �1��g��  2�V�z���?�c�
/��VISBCK������*.VD/[/��FR:\F/�.��Vision� VD file �/��/�/�?�)? �/:?_?�/�??�?�? H?�?l?O�?�?7O�? [OmO(O�O O�ODO�O �OzO_�O3_E_�Oi_ �O�__._�_R_�_�_ �_o�_Ao�_Rowoo �o*o�o�o`o�o�o�o�oO��MR_G�RP 1G���L4uC4  B�8p	 ����|�p�۬B��D���fnӺ�MT� ��� ����u�y�q� ��r�x%��tA�5s�s�_�J�N��L��K�~M��&�H>;�E���L������p@4���B��A�z�?�Bf���9�f���A��%�A�A��A��A������F�@ %���-��g��fF6�D�M�qD�� BT�_�@��Ý�?@��u�Ï6��؝����5��5�����Ɵ��ß��� ��A�?�M���r����������  �@���@h0�?�\	@�B� ɯ�����8�#�\�G� ��k�������ڿ���v4uBH8p 9���:�L�^���̲Z�?�W[�`�w�̉�;�A@O���@��33@����\����ɿ�Ɋ��"� ��I�[�F��jߣߎ���߲�<�G�=��<�m]<��+=~�m<�c^��8eN7���7ѷ7ߑx7;�51����:���7�p��t2��pY�p��p�O��RO��w�⮓p �p5O�0'���t� ��-���C��#� 1���Y���������� ����0T?xc ������� >)bM�N�P� ^�Z��/�+/ /(/a/L/�/p/�/�/ �/�/�/?�/'??K? X9�X?~?�?�?i��? �?=?�?�?OOBOTO ;OxOcO�O�O�O�O�O �O�O__>_)_b_M_ �_q_�_�_�_�_�_o o��7o�{�%�7��o [��o��o�_ �o$ H3X~i�� �������D� /�h�S���w������ ㏩�
���.��R�=� v�a�s�����П���� ߟ��(�N�9�r�]� ��]?��̯ޯ�?� {�$�J�5�n�U���y� ��ȿ���׿���4� �D�j�Uώ�yϲϝ� ����������0��T� o-o��Qo��uo�o�� �o��o5�G�P�;�t� _����������� ��:�%�^�I���m� ��������� Ǐ! �ZE~i�� ����� D /hS�w��� ���
//./@/�d/ ��/s/�/�/�/�/�/ ?�/?<?'?`?K?�? o?�?�?�?�?�?O�? &OOJO5OnOYOkO�O k�}��O���O����1_ ��U_�O�_y_�_�_ �_�_�_o�_0oo@o foQo�ouo�o�o�o�o �o�o�o,Pq ;�[����� ��:�%�^�I�[��� �����܏Ǐ ��� 6��Z�l�~�E/O��� �؟ß�����2�� V�A�z�e�w�����ԯ �������,�R�=� v�a������������ �O�O'�I_K�_7_9_ ?ϥ�o_տ������� ��8�#�\�G߀�kߤ� �ߴ���������"�� F�1�j�U�g��g�� ��������B�-� f�Q���u��������� ����,P;t �M������� k(L3\�i �������$/ /H/3/l/W/�/{/�/ �/�/�/�/?�/2?D? �e?/ϩϛ?eϿ?�� �?��
O%?.OORO=O vOaOsO�O�O�O�O�O �O__(_N_9_r_]_ �_�_�_�_�_�_��o �_8o�_\oGo�oko�o �o�o�o�o�o�o" F1C|g��� ������B�� ;�x�c�������ҏ�� �����>�)�b�M� _�����������˟� ��:�%�^�I���I? [?��?ٯ�?�?��? 3��?Z�u�~�i����� ƿ���տ� ��D� /�h�Sό�wϜ��ϭ� ����
���.��_oo '߈�s߬ߗ��߻��� ���*��N�9�r�]� ����������� �8�J�\�n�5����� ������������  F1jU�y�� ����0T ?xc��������$FNO �������
F0! �  T�1 D|����RM_CHK�TYP  ��\������!{OM _MIN" ��N �  �X�SSB_C�FG H� ��{/���r#�/�/�TP_D�EF_OW  �-"�(IRCO�M! �/�$GENOVRD_DOC&s�ѡ<THRC&� d5d4_EN�B�/ 0RAV�C_GRP 1Id'�! X��?� �?�?�?�?�?O&OO JO1OnOUOgO�O�O�O �O�O�O�O"_	_F_X_ ?_|_c_�_�_�_�_�_��_�_�_0o2ROUrp0O�Q ������"��8��?T��o3o|o�o�o 7 D��`3�1�o�v/��@r�|B��ҡrĩoi4og0SMUTm3Pt=���������|�$HOS�TC]"1QOip [��o 	�x�{��0�'�O�eC�t���������b��ۏ����4�5�Ȁ	�anonymous8�f�x�������� ���.�P�ʏ7�I� [�m���������ǯٯ ��:�L�!�3�E�W�i� ��ʟܟ���տ$��� ��/�~�@�e�wω� �Ͼ���������� +�z�����D߲ϗ�� ����������'�9� K�]�߁��ϥ���� ����<�N�`�r�t�Y� ��}������������ ��B�0��gy ������"�4�6 j�?Qcu��� �����T)/ ;/M/_/q/���� ��/,??%?7?I? �m??�?�?�?�// (/�?O!O3O�/�/�/ �/�?�O�/�O�O�O�O _Z?/_A_S_e_w_�O �?�?�_�_�_�_j}�q�ENT 1ROk� P!�_Eo  @p3opo_o�oWo�o {o�o�o�o�o6�o Z~A�e�� ��� ��D��h� +�=���a���揩� 
�͏�@�/�d�'��� K���o�������ɟ *��N��r�5���Y��k�̯��𯳯�ת?QUICC0!����p�3�1q�M�_����3�2�������!?ROUTER�����`�!PCJO�Ga�<�!19�2.168.0.�10:�gNAME� !"j!RO�BOT��nS_C�FG 1Q"i ��Aut�o-starte�d`DFTPkO HтO�_s߸O�ߩ߻� ����$_��'�9�\� J��߁������JF !�3�E��Y�{�1�b� t�����g�������� '���:L^p� �QOcOuO� O� $6HZ)~�� ���k�/ /2/ D/V/����/��/ �/�/
??��/R? d?v?�?�/�???�?�? �?OOg/y/�/1O�? �O�/�O�O�O�O�O�? _&_8_J_mOn__�_ �_�_�_�_)O;OMO_O a_Fo�Ojo|o�o�o�o �_�o�o�o/o�o�o Tfx���_�_o !o#�Wo,�>�P�b� t�C������Ώ��� ���(�:�L�^��� ���ʟ�� �� $�6��Z�l�~����� şG�د���� ����T_ERR S���.�>�PDUSI�Z  �^���U�>n�WRD �?ը��  �guest \�����ҿ���Ͽ��SCD_GROU�P 2TM� ����1�!��L9_N��  ��>R�	 i-	��v�����E E�ATSWILIB���\�N�ST �4�@��bǀ�}�FRS:�T�TP_AUTH �1U=�<!iPendan�޶�����!KAR�EL:*�(�:��KCO�_�q�G�V�ISION SE!T8��ߦ��!���� ��D�"��:�4��X��j������CTR/L VM�����
��FFF�9E3�璉��D�EFAULT-��FANUC W�eb Server-�
�Ė�����������������<�WR�_CONFIG �W�����-�>�IDL_CP�U_PCL���B�ȩ�g �BHMM�INXE�lGNR_IOG�|���S�O �NPT_SIM_�DO��TPM�ODNTOL� >�_PRTY�g�KOLNK 1XM�	�-?Qcu���MASTEҜ ���	O��O_gCFG��UO��|��CYCLE���F�_ASG 19Y*�
 �\/ n/�/�/�/�/�/�/�/��/?"?4?F?�/"N�UM{�Q�{��I�PCH/���RTRY_CNL�Q���SCRN_UP)D{�,�U� ����ZM�r�O����$J23_DS/P_EN��M���~@OBPROC$C���JOG4�1[�M� @��d8��?�Q;�OQ??>ZCPOSREDO��KANJI_�K���CM��3\*�x�E�O�ECL_Lw �l2�?�@EYLOGWGIN����|A�U��$LANG?UAGE ��g�F� �Q>�LG��2]�ﱢ����xRBа���Pm ����'0�H���0��MC:\RSCH�\00\.��PN_DISP ^M�॔��|�z�<�LOC��^Dz�=#��{�iPBOOK  a�>'}@���������`XJi�o�o�o�1~D}7xVy�	�e�i��Me��}b�G_BUFF 1-`�2��� �b�����'�T�K� ]�����������ɏ�� ����#�P�G�Y����)d`@DCS b>�m =���S|�������� �8C��I�O 1c:+ 	O]����]�m���� ����ǯٯ����!� 5�E�W�i�}�������@ſտ����8�E� _TM  9kdC� Y�k�}Ϗϡϳ����� ������1�C�U�g� yߋߝ߯����߾t=��SEV�09m7�TYPC�U�6�H�Z��}�ARS| R_�s�2�FL 1dF��0�Ο��������(�L:�k�TPfPC�%�}rmNGNAM$D�e	��UPS1`G�I�5 Q�5��_L�OADA@G %�9j%CAL_T�C���D
MAXUALRMl7�z8 ����3�0�Tq C4ae��i�~S tb@g@f:+ �w	%�����- Q<uXj�� ���/�)//M/ 0/B/�/n/�/�/�/�/ �/?�/%???[?F? ?j?�?�?�?�?�?�? �?�?3OOWOBO{O�O pO�O�O�O�O�O_�O /__S_e_H_�_t_�_ �_�_�_�_o�_+o=o  oaoLo�ohozo�o�o �o�o�o9$]�D_LDXDI�SA��E�6�MEM�O_AP��E ?=��
 �fy ������&�8�~ ISC 1g�� �P��Lt���� ��O؏Ï��� �2� ��A��z�e������� ԟU�㟷��.��R� 9�v�������k�Я�� ��ۯ�*���9��r� ]�������̿M�ۿ�� �&��J�1�n��}� ��c��ϳ������"� ��1��j�Uߎߠ�Y��_MSTR h��ݳ�SCD 1i�}�����&��J� 5�n�Y�k������ ������� �F�1�j� U���y����������� ��0T?xc ������� >);t_�� �����//:/ %/^/I/�/m/�/�/�/ �/�/ ?�/$??H?3? X?~?i?�?�?�?�?�?��?O��MKCFG� j��O��L_TARM_5Bk��wKB C��p�NxpMETPU܅pB����NDSP_CMNT�EpI@CF�E�� l�ނ�NBKA_T�EP�OSCF�G�NP�RPM�O�HPST�OL 1mc�4@@<#�
�Q	A�U �_�W�_�_�_�_o�_ �_<oo0oroTofo�o �o�o�o�o�o�a�A�SING_CHK�  \_$MODAQhCn;O�GKJNu�DEV 	��	�MC:~|HSI�ZE�@���NuTA�SK %��%$�12345678�9 ��uLwTRIoG 1o�� �F3%��OL�  1�r�U����vYP�q]����MsEM_INF� 1poG �`)AT&�FV0E0���)�ށE0V1&A�3&B1&D2&�S0&C1S0=>�)ATZ��J�1�HN�v��j���-�A��Ο���ٟ�(� ܏M� ��$�6��� Z�˯�����%�� I�[�B��2�D���h� z������¯3�j�W� ����HϱϘ����� ��߾�п���e�� ���Ϛ߿�r��ߞ�� � �=����s�&�8� J߻������(���� ��K��o�V�����X� ��|����#��G Y��}0��\�����#NONITO�R�@G ?�{  � 	EXEC�1C>2D3D4�D5D�F7D8
D9C?��C �O�[�g�s ���������2�2�2�2��2�2�2�2�(2(2(3�3�3ONqR_GRP_SV 1qˉ�,�(q>�9�?��h���?���<��@�g,Ѯy}�q_D���~0APL_NAM�E !�E;0��!Defaul�t Person�ality (f�rom FD) �-DRR2�! 1r�)deX)dh�;1�AX dO�?�? �?�?�?�?OO%O7O IO[OmOO�O�O�O�O�O�O�O	X2�?-_?_ Q_c_u_�_�_�_�_�_=r<_�_oo/oAo Soeowo�o�o�o�o}x�R�" 1w39jp=\@r0 ���@r��a @D�  &q?�s�a?@pq�@qAI�Ez � 3qqEw;�	l~'r	 0Ap�er@es_qp�{t��{t� Ki�K��J���J����J�4�J~���Ezvq�^q�P���|�p@�z��r�f�@�S���/q��s�=�N���
������T;f�
�����p�*  �_p  �U�>Q���U���?��?�����OO�����R�����(q����Buʍ�|}  ����pj  T�������܏ 	�'� � C��I� �  {��ߍ:�Èg�?È=�����r@�����~q��D*�rÈ��~N_0�  ''��q(��@a�@�t�E@4�@8���pCP�KCa�fa�\�B`��Cd�p�@�V��voo$~�}����wAAV���_0ϡ*��pp�qD8u�����5� �Y��}�� ��t O� �ru �4 ������Ӄ� �::u�qp�p �?�ff Q��Ŀֿh� ������q�4�B�>������yPplϖ���xvqevم�>L������r<	�I<�g�<#�
<2���<D��<���
����s��s_��?fff?榐?&��t@T���/�?�`?U?ȩ?X�?��� ���(tk�ts�w�� �[t���߲������ ��3��W�i�T���\�F_0|���x����d������A���G�@ G��F���� t������������� +�z��O�  ڏ��(��d' 9K��`r��P����Ϣ�$ ��&/w�M/�q/\,�w��z/�/�/�/�)�2V��$-�pB�a�01?m��"�� �!71�@I�;M`B�@��@`�9�@y��?�h�? �@�3��[N��N�N�E��<�/k?�}0�>��ڟ��A�p�C�F�@�S��?u�X������@�t��%�h�?�K�G��Gk�nF&�Fצ�pE,8{�? �F�ZG����F�nE�D�E,ڏO@����G��F7���F��ED�� _��/tO_O�O�O�O�O �O�O�O__:_%_J_ p_[_�__�_�_�_�_  o�_�_6o!oZoEo~o io�o�o�o�o�o�o�o  D/hSe� �����
��� @�+�d�O���s����� Џ��͏��*��N� 9�r�]�������̟�� �۟���8�#�5�n��Y���}�����گŮ(��13�jiꯣ��y��ӥ3Ա��<��4 ��7�I���P�c�u�W��jb����1w�����������@���C�1̤P��	PuΔ����� ������#�М��� >�)�A�M�_�5$x�B� �߮��������ņ ��{�5�C�U�y_�q� �������e����-��Q�?�u�_�2v�0�$��G��ߢ� B !!� B
�CH � K���� &8J���~@������$��E� � �ў�c�%
 �0BT fx��������//�:
 ���o�x}��$M�SKCFMAP � ���� ��
��-S#ONREL  g��j!��S"EXC/FENB�'
h#�%ε!FNC�/�$JO�GOVLIM�'dt� �"dS"KEY�'u5S"RUN�,�5S"SFSP�DTY���&�%�#S�IGN�/�$T1M�OT�/�!S"_C�E_GRP 1x��j#\ϯ�?ǯ OOe�??O�?cOO XO�OPO�OtO�O�O�O _)_�OM__q_�_:_ �_^_�_�_�_oo�_ 7o�_[omoTo�o^S �TCOM_CFG 1y`-�o�o��o
�a_ARC_�"g��)UAP_�CPL�$NOCHECK ?`+ f�lxj| ����������0�B�T�f�x��+N�O_WAIT_L�w7f%�2NT�az�`+ʁ_ERRr�2{`)��� �o#�5�G�S�9#k�}�^ItT_MO��|��,  &ށoȟ��_PARAM�2}`+�	���~g���E� =��345678901_�q��� Z������������د0 �2��}g�d�v��	���JsUM_RSPACE]/ӿݴ��$ODRDSP�sz6�(OFFSE?T_CART9��DIS��PEN_FILE<�z1�a���pOPTION�_IO?�PWO_RK ~�7�# �Э�t��
g�8������	 ������t����RG_D?SBL  ��#�6��RIEN�TTO� ��C��i!=#�p�UT�_SIM_D{��g":"�V��LCT ԍ�����a��>��_PEXE=���RAT���&�%M0��>�UP ������%�7��[�i���$�2�3r)d�eX)dh���X d�������� ����
��.�@�R�d� v���������������$2��HZl ~��������<7&8J\n �������'���0O�1w(��O�(�_Ҙ��20 �Ԧ  � @D�  .!?��4#!?��6!��D4  EzP#Ijd,�;�	lF"	 '0��"@�#~!�* ��$��$1�H)�!H,�H�8�Hm�G�?	{G�8�$�g��~f��/ <1�C�Z�1�Z�� 3N!-?���*  �p � �L0>H0� # �+=C?U2�]��-�B]�Btr�«{���¼�2?�?�2G!�31�])�a/1�@�  �@��j  K0�&F��DO~e	'� � bB�I� �  ����==���8�O�K`�@�O�@ �>��OIK�0�N�&ykN ._4Q'~�HT,1o0CZ�fZ�S0BW0*>S_eR\�IJ�a��@uA�&o�o$�-���{gAu@�Z5P�QIJ �AeJ" W%3O0ooTo?oxocm��� �t �O� ru �4 ��b<�e��� :�5�����0 �?�fAf�qk�o�o�o�ʈ3��Q8��Saz>��`�agiP����g�Q�!�&�5�>L��@�32<	�I<�g�<f�<2���<D��<��`���/�5"��|~r`?fff?�@�?&<�kd@T��N�?�`?U��?X�^���R 7�G$fi6%��4'�� � z$�я
���.�� R�=�v���s������� �͟�}�������`�~��G�@ G�0 ��������ί���� �(��L�7��Rn�1� _��?��?#��G�� ��4�F�X�j�	�ϑπ+��ϯ���������R�4��TEߖ��l�xߐ�{�?�ؙ�P���������uD�C��1��P'�&�1�ظ���в�V�@I��Z�M`B@���@`�9@y���?�h:� ��@�3�[N���N�N�E��<��/����>���ڟ�A�p��C�F@�S����8�X������@�t��%��h�°�1G���GknF&��FצpE,8�{� F�Z�G���F�n�E�DE,ڏ�*�<��G���F7��F��ED��~v�ߓ�~� ������������5  YDi�z�� ����
U @yd����� ��//?/*/c/N/ �/r/�/�/�/�/�/? �/)??9?_?J?�?n? �?�?�?�?�?�?�?%O OIO4OmOXO�O|O�O �O�O�O�O_�O3__ W_B_T_�_x_�_�_�_��_�_�^(��3�j�i	o�q��:e�U3�Ա�*o<o�q4 ��Voho�q�Pqło�ovbjb�o��o1w������m�i>,b�P|õP�rP�~�� ���o��o��Bi#���$�]�H�`�l� ~�Tԗ�aߏ͏�� '�=i�u������T�b�t�y~���Ɵ��ʟ؟ ꟬r���2�L�:�p�h^���~z2��$�f'G����`B?�3��B)�CH4��`j� ��+�=�O�a�s�ɳ��������ӿ���*�d��`�`��r�����e
 �� O�a�sυϗϩϻ��� ������'�9߸�)�� ����x}���$PARAM_MENU ?���  �DEFPU�LSEE�	WAITTMOUT���RCV�� �SHELL_WR�K.$CUR_S�TYL����OsPT���PTB���C��R_DECSN�ЅuX�R�d�v� �������������/�*�<�N�w�r�US�E_PROG �%��%s�����CC�R���u����_H�OST !��!����T�p��)���+e��_T�IME��1��  �r�GDEBUG�/ �ۇ�GINP_�FLMSK��	T�R��PGA�  2����CH���TYPE~��� r�l������� � //;/6/H/Z/�/ ~/�/�/�/�/�/�/? ? ?2?[?V?h?z?�? �?�?�?�?�?�?
O3O��WORD ?	>	RS� �S/PNS�U��oBsJO��RTEL �0TRACECToL 1����� �p ��p�p�N�FDT� Q���@�@�D(���P�R6��smU�q-P )�3R%�WP0RP8R�P@RP�R�R�	T	T		T	T*	T	T	T	T1 �R	T	T	T�	T	T	T	T�	T	T=�R	T�	T�R!	T"	T#�	T��R&	T''� E_W_i_{_�_�_�_�_��_�_�_oo/o	T%TIhQ(	T)	T*	TU+	T,	T-	T.	T/	T0Qocouo�o�o �o�o�o�o�o) ;M_q���rQU1	T2	T4	T5	TU6	T7	T9	T:	TU;	T<	T=	T>	T%?	T@	TY�� ����!�3�E�W� i�{�������ÏՏ� ����/�A�S�e�Q ]Q�c�u��������� Ͽ����)�;�M� _�qσϕϧϹ����� ����%�7�I�[�m� ߑߣߵ��������� �!�3�E�W�i�{�� ������������� /�A�S�e�w������� ��������+= Oas����� ��'9K] oE������� �/#/5/G/Y/k/}/ �/�/�/�/�/�/�/? ?1?C?U?g?y?�?�? �?�?�?�?�?	OO-O ?OQOcOuO�O�O�O�O �O�O�O__)_;_M_ __q_�_�_�_�_�_�_ �_oo%o7oIo[omo o�o�o�o�o�o�o�o !3EWi{� �������� /�A�S�e�w������� ��я�����+�=� O�a�s���������͟ ߟ���'�9�K�]� o���������ɯۯ� ���#�5�G�Y�k�}� ������ſ׿���� �1�C�U�g�yϋϝ� ����������	��-� ?�Q�c�u߇ߙ߽߫�����������$PG�TRACELEN�  ��  �_������_UP �����@�H�,��A��_CFG M�@�*���A��m�#� m����m�U�DEFSPD� �`��q#����INX�TRLW �`���8}����IPE_CON�FI\��@���@�m���LI�DY�`�<�GR�P 1��*�����@�
=�[����A?C�C�
�XC)��Bg����#�����d}����/�/�� 	 ��������� ´����B  8N8r���> �6>7��D���� ='?�=)��� �O:s^���~���  Dz#/��
/G/� W/}/h/�/�/�/�/�/ �/?�/
?C?.?g?R?��?��
V7.1�0beta1m���0B=q�2`�ff@��2>�{���1=����1�A>ff�1@�f�f�2�\)�2D�_�?�  A@	AL�0�1Ap�3�ș?`7OIO[OmO|K�����,��?�O|?�O�O _ _9_$_6_o_Z_�_ ~_�_�_�_�_�_o�_ 5o oYoDo}oho�o�o �o�o�o�o&/1�o U@R�v��� ����-��Q�<��u����?�3F@  ��������@��M� �0�&�N�`��O�O�O ������ޟɟ��&� �J�5�G���k����� ȯ���ׯ�"��F� 1�j�U���y������� ���ͿB�-�f� Q�cϜχ��ϫ����� ���,�>�)�bߍ��� я�߭������� A�:�e�w�������C� ������������6� !�Z�E�W���{����� �������� 2V Aze������ �
�.R=v as������ //</N/yߋ߽߇/ �/���߻/�/�/-�&? Q�c�u��?//�?�? �?�?�?�?�?"OOFO 1OjOUOgO�O�O�O�O �O�O_�O0_B_-_f_ Q_�_u_�_�_��_�_ �_oo>o)oboMo�o qo�o�o�o�o�o�o (S/e/w/�/s�/�/ �/?�? ��=?O? a?s?l���{����� ؏�Տ���2��V� A�z�e�w�����ԟ�� �����@�R�=�v� a����_��Я���� �*��N�9�r�]��� ����̿���ۿ�? Qc�_ϙ���� �������)�;�M�� X��|�gߠߋ��߯� �������	�B�-�f� Q��u��������� ���,��P�b�M��� ������k����� :%^I�m� ���� +�=�O� 9K�ϗϩϟ��� ���'�9�2/�// h/S/�/w/�/�/�/�/ �/
?�/.??R?=?v? a?�?�?�?�?�?�?�? OO<O'O`OrO���O �OWO�O�O�O�O_&_ _J_5_n_Y_�_}_�_ �_�_�_)[%o7o�q���o�o��$�PLID_KNO�W_M  ����Q�dSoV ���`��O! 3�_WBT��R-��cM_GRP 1���j& dzp��oo$tv�t_���d��d M`�z	�}{�v,�S��e �o�C�?���c���ۏ �������5��h�e� )�K���u��������� ���+���g�;���`I�[���Ӯ�aMR�sŎ�}T�Uxa|O  xb3�E�Y�T�*���N� `�r��������̿.� @�U�P�&ψ�J�\�n� ���ϼ϶���*�<�Q�`L�"߄�F��ST�q�1 1�����v�`0� @��� �U�������H�+�=� ~�a�s�������� �����'�h�K�]������2�����Q�<����3����������4/A��A5Zl~���6������7�
.��8GYk}�ӿMAD  $��� ��PARNU/M  ��|����SCH� �
�<'!J)�c\%UPD�/%�q�/�$��_C�MP_�p�m`�'��e�$ER_CHK�%���j�"�/��+RS��o�a_M�O�.?@5_*?�__RES_G�А�� */���?�?�?�?O �?%OO*O[ONOOrO@�O�O�O{7���<�? �O}5
 �O__3Y  &_E_J_3� e_�_�_ 3� �_�_�_3F�_ oo3�"oAoFo2�V 1��e�q"@�cX��`P�`�`W���`l�` @cV���`�@2THR_�INR���rr5d��fMASS�o Z��gMN�osMON�_QUEUE Q��u�&�p��p�N� U1N v�+cp�ENDeqg?yEX1E�u� BE�po>`sOPTIOlwp;�cpPROGRAM7 %Cz%bp�o�+/arTASK_I���~OCFG �C/7�j�DATuA���s�@��2�������'�я J�\�n���+�����ȟxڟ쟟�INFO������Rt��@�R�d� v���������Я��� ��*�<�N�`�r���Ж�������� ��Ii�� DIT �s�ϛ�WERF�L�x�c��RGAD�J ���A�  ]�?v�i��aA�cq�n����'�?���v�<��/�%���5ȲO��±��2���!�t 	 h���b�����Ard�t$B�v��*U�/W� **�:`�P�bր�;����ҍ՝߉5��NӼ� ���ߕ��������� ��A�7�I�[���� �������=�����v� !�3���W�i�{����� ��������o� ASЇ�� � �C�'I��U�y��RIORITY� w�&�E�MPDSP�q3ϱUw-��;OG�_TG0�W��Gz�TOEp1���� (!AF��`Ef09/D'!�tcpD/l-!�ud[/�.!iccm�/�o�XY��������)� 0m��/
?����/3? 5"?_?F?�?j?|?�? �?�?�?OO�?7OO�[OmO*D�PORTT�q���%E��_CARTREP��p���aSKSTA�x�zSSAV?p����	2500H809�(����D������`.�kY_xk_i�PURGE�p�B0��yWF�PDOU���W2 �T��J�WRUP_DEL�AY ����TR_HOT��b��8o��UR_NORMA�L�(o}oLfSEM�I[o�o�oqQSK�IP���� x kg);M} ~l������ � �2�D�
�h�V��� ����v����ԏ
�� .��R�@�b������� r�П������ޟ(��N�<�r�������$�RBTIF���R�CVTM�$����DCRƳ��l��qB
�B}��>A��@��_��"���x��$��Q�V����HU���o���6�`�\ �<	�I<g��<#�
<2���<D��<���
r�Y�¿Կ  ֿ��� �2�D�V� h�zόϞϰ��ϭ��� ��
����@�+�d�G� �ߚ�ݿ��������� �*�<�N�`�r��� �ߺ���������� 8��\�n��ߒ����� ��������"4F XC�U��y��� ���0B��f x������� //,/P/;/M/�/ q/�/�/�/�/�/?G Y:?L?^?p?�?�?�? �?�?�?�? O�/$OO HO3OEO~OiO�O�O�O �O?�O_ _2_D_V_ h_z_�_�_�_�_�_�O �_�_oo@o+o=ovo Yo�o�o�O�o�o�o *<N`r�� ��o������ 8�J�-�n����o���� ȏڏ����"�4�F��X�j�y��GN_A�TC 1��� �AT&FV�0E0y�AT�DP/6/9/2{/9��ATAy��,AT%G�1%B960���+++ޟ,ّH��,�IO_TY�PE  \�ƣ�e�{�REFPOS�1 1�G� O x�f���_� Ư[���������B� -�f����%���I���俒�����ҿ3�� W��{�ϟ�:Ϝ��� p��ϔ�߸�A�����  �:ߛ߆߿�Z���~� ���=���a��߅�  ��D�V�h����� '���K���o�
�l��� @���d��������� ��
kV�*�N �r��1�U �y&8r�� ��/�?/�</u/ /�/4/�/X/�/|/�/ �/�/;?&?_?�/�?? �?B?�?�?x?O�?%O �?IO�?�?OBO�O�O �ObO�O�O_�O_E_ �Oi__�_(_�_L_^_ p_�_o�_/o�_So�_ wooto�oHo�olo�o �o�o�o�os^ �2�V�z�� �9��]����g�y�2 1���.�@�z� ����"�@�ۏd��� a���5���Y��}�� ����ş��`�K���� ��C�̯g�ɯ���&� ��J��n�	��-�g� ȿ��쿇�ϫ�4�Ͽ 1�j�ώ�)ϲ�M��� qσϕ���0��T��� x�ߜ�7ߙ���m��� ����>�������7� ����W���{���� �:���^������� A�S�e��� ��$�� H��li�=� a����� hS�'�K�o �
/�./�R/�v/ /#/5/o/�/�/�/�/ ?�/<?�/9?r??�? 1?�?U?�?y?�?�?�? 8O#O\O�?�OO�O?O �O�OuO�O�O"_�OF_ �O�O_?_�_�_�___ �_�_o�_	oBo�_fo�o�o%o�o����3 1���[omo�o% IOom�,�� b����3��� �,���x���L�Տp� ������/�ʏS��w� ���6�H�Z������� ���=�؟a���^��� 2���V�߯z������ ¯��]�H������@� ɿd�ƿ����#Ͼ�G� �k���*�d��ϰ� �τ�ߨ�1���.�g� ߋ�&߯�J���n߀� ����-��Q���u�� ��4����j����� ��;�������4����� ��T���x�����7 ��[���>P b���!�E� if�:�^� �/���/e/P/ �/$/�/H/�/l/�/? �/+?�/O?�/s?? ? 2?l?�?�?�?�?O�? 9O�?6OoO
O�O.O�O�RO�O�o�d4 1� �o�O�O�OR_=_v_|O �_5_�_Y_�_�_�_o �_<o�_`o�_ooYo �o�o�oyo�o&�o #\�o��?� cu��"��F�� j����)���ď_�� �����0�ˏݏ�)� ��u���I�ҟm����� �,�ǟP��t���� 3�E�W����ݯ��� :�կ^���[���/��� S�ܿw� ϛ������� Z�E�~�Ϣ�=���a� ���ϗ� ߻�D���h� ��'�a��߭��߁� 
��.���+�d��߈� #��G���k�}���� *��N���r����1� ����g�������8 ������1�}�Q �u���4�X �|�;M_� ��/�B/�f// c/�/7/�/[/�//?<�O T5 1�_�/ �/??j?�?�/�?b? �?�?�?!O�?EO�?iO O�O(O:OLO�O�O�O _�O/_�OS_�OP_�_ $_�_H_�_l_�_�_�_ �_�_Oo:osoo�o2o �oVo�o�o�o�o9 �o]�o
V�� �v��#�� �Y� �}����<�ŏ`�r� �����
�C�ޏg�� ��&�����\�埀�	� ��-�ȟڟ�&���r� ��F�ϯj�󯎯�)� įM��q����0�B� T����ڿϮ�7�ҿ [���Xϑ�,ϵ�P��� t��ϘϪϼ���W�B� {�ߟ�:���^����� ����A���e� �� $�^�����~���� +���(�a���� ��� D���h�z�����' K��o
�.�� d���5?-46 1�8?��. ������/� /N/�r//�/1/�/ U/g/y/�/?�/8?�/ \?�/�??}?�?Q?�? u?�?�?"O�?�?�?O |OgO�O;O�O_O�O�O �O_�OB_�Of__�_ %_7_I_�_�_�_o�_ ,o�_Po�_Mo�o!o�o Eo�oio�o�o�o�o�o L7p�/�S �����6��Z� ���S�����؏s� ���� ����V��z� ���9�]�o����� ��@�۟d�����#� ����Y��}����*� ůׯ�#���o���C� ̿g�𿋿�&���J� �n�	ϒ�-�?�Qϋ� ����߫�4���X��� Uߎ�)߲�M���q��� �ߧ߹���T�?�x�� ��7���[���������>���b�HZ7 1�e�!�[����� ���!��E��B{ �:�^��� ��A,e �$ �H��~/�+/ �O/��/H/�/�/ �/h/�/�/?�/?K? �/o?
?�?.?�?R?d? v?�?O�?5O�?YO�? }OOzO�ONO�OrO�O �O_�O�O�O_y_d_ �_8_�_\_�_�_�_o �_?o�_co�_�o"o4o Fo�o�o�o�o)�o M�oJ��B� f�����I�4� m����,���P���� �����3�ΏW��� �P�����՟p����� ����S��w���� 6���Z�l�~����� =�دa����� ����� V�߿z�Ϟ�'�¿Կ � ρ�lϥ�@���d� �ψ���#߾�G���k��ߏ�u���8 1� ��<�N߈����*�0� N���r��o��C��� g������������ n�Y���-���Q���u� ����4��X��| );u���� �B�?x� 7�[���� >/)/b/��/!/�/E/ �/�/{/?�/(?�/L? �/�/?E?�?�?�?e? �?�?O�?OHO�?lO O�O+O�OOOaOsO�O _�O2_�OV_�Oz__ w_�_K_�_o_�_�_o �_�_�_ovoao�o5o �oYo�o}o�o�o< �o`�o�1C} ����&��J�� G������?�ȏc�� �������F�1�j�� ��)���M���蟃�� ��0�˟T����M� ����үm�������� �P��t����3�����ߴ�MASK 1����� ���?XNO  ��~�MOTE  /�����e�_CFG ��lͷ���PL_RANGh�b�p��POWER �����x�SM_D�RYPRG %�l�%i����TAR�T ����UME_PRO�� �{����_EXEC_E_NB  `�tɏGSPDTЖО����TDB����R�M����MT_�T���j��OBOT�_NAME �l�j�׹OB_O�RD_NUM ?����=�H809  `����	d�H	��\췰���� ,��:��	@���D|����PC_TIMoEOUT�� x�oS232��1�0���� LTE�ACH PEND�AN������)��[�R� M�aintenance Consb��&�_�"B�T�KOCL/C.Д�r��5��� No Use��r���]���NPO������v���CH_�LW��lβ�	�a0MAVAIL�w�����t���PACE1 2�l� +���	������p�8�?��,	;, q�i���� �	�-OA/b/%/ ��/)0�4��-�� �	/{/-/O/A?b?%?@�/�??�?:�2���/�/?�?+?M? \O}O@O�O�O�O�O�;3�?�? OO$O�OHO jOy_�_]_�_�_�_�_�;4�O__/_A_�_ e_�_�o�ozo�o�o�o�;5o(o:oLo^o �o�o����
����;63EWi {)���Џ񏴏�'��<��;7P�b�t� ����F���ޏ��џ #�D�+�Y��;8m�� ������c�ٟ��
�+���@�a�H�v��;h �Nl� m��
Ӱ ¿����� %�7�I�[Ϲ(˧~ͱ� ����S����d��ؿ ��*�<�N�`�r߄� zόϞη/�ߓ����� �0�B�T�f�x��� �߼���������� "�P�b�t������������������
� `n� @�S�� a=�E��!*� ����
��)G �/q�MWi� �����7/I/g/ /O/�/�/m/w/�/�/��/�/��
�R?�;_MODE  ��^h9S ���A?����ޯ}�?�?J�	OAO�DCWOR�K_ADx=	5���AR  ��𚠏@FOy@_INT�VALx0����:R_OPTION�F� �5`V_D�ATA_GRP �2�����D9�P .O_*O>_)Y+?k_Y_ �_}_�_�_�_�_�_�_ �_1ooUoCoyogo�o �o�o�o�o�o�o	 ?-OQc��� ������;�)� _�M���q��������� ˏ��%��I�7�m� [�}�����ǟ���ٟ ����!�3�i�W��� {�����կï�����/�1�$SCAN�_TIMw1I��5�I�R �(�3�0(�L8�ѰѲ�34Q	���1���:�3_�����?��Ӳ2Ĉ���d����/R�� @���Q�c�u�RU0�D� �P��0[ � 8�@��������D�����+�=�O� a�s߅ߗߩ߻��ߒ��1B����#����S����;��oRT���1p���?t��DiD��>��  � lӲ�1 �񘱐����������� ���#�5�G�Y�k�}� �������������� 1<��Sew� ������ +=Oas��� ���>P�� /2/ D/V/h/z/�/�/�/�/ �/�/�/
??.?@?R?�d?v?�?�?�5�?  0�2'���?�?O#O 5OGOYOkO}O�O�O�O �O�O�O�O__1_C_ U_g_��_�_�_�_�_ �_�_	oo-o?oQoco uo�o�o�o�o�o�o�o v_�_/\n� �������� "�4�F�X�j�|�����`��ď֏�7�?  � 
��.�@�R�d�n��� ������ɟ۟�����#�5�G�Y�k�}��� 葯�è�ί�� ��(�:�L�^�p����ɶ����¿������ ����	�12345678����������02�D�V�h�z��������������� ��0�B�T�f߭��� �߮����������� ,�>�P��t���� ����������(�:� i�^�p����������� ���� A�6HZ l~������ �+ 2DVhz ������
/ /./@/R/d/v/�/�/ �/�/��/�/??*? <?N?`?r?�?�?�?�����?�?�3�/OO�)OMyCz  B}p��   �Qx�2���:�$SCR�_GRP 1�(��e@(�l��0�@} � ۱��	 �C�A�B�D�1����I���F�O�O$_I}[���C�PP�������fX![w\L�R Mate 2�00iC �90���U�LR2CA ���C���
�X��S�AշV�wS��!Q�J�Ai	�RLo^opo�o�o�lް��@5n߲�o �O!_
�G�?���@`�o�=Hv?Fh�-,�IB�K@���r��t�AA\@�  @����A@WP�  ?~�6��rHK@G��z��AF@ F�` q�y�p��������я �����?��}�>�`j�U�g�y���B��� .�ߟʟ��'��$� ]�H���l�����ɯX^�ū��_�����e
��Y��6�@��=�ò"`��G"���B�6���90��>G��@EL_DEFA�ULT  �d�_�/�ޱ�MIPOWERFL  �E��ݲ�oWFDO� ����AERVENT �1����`����0L!DUM_�EIP��p��j!AF_INE�<���!FTdϽ������!�o� ����-�!RPC�_MAIN.�غ8�y�@�VISI��y�h���!TP�ГPU��w�d���!�
PMON_PR'OXY�z�e �]����+�s�fL��!RDM_SRV��rw�g����!RҸd�|�h��A�!
B��Mt�t�i0���!?RLSYNC�����8|���!ROSc� �4��%�� I��(r�^� ����'�  o6HZ������/�5/;�ICE_KL ?%K�� (%SVCPRG1:/�*l%lCD�/�-3�/�/q 4�/D�/q 5�/�/q 6"?'?q 7J?O?q �T�?�,9�?�;n$��? q!t/�?q!�/Oq!�/ ?Oq!�/gOq!?�Oq! <?�Oq!d?�Oq!�?_ q!�?/_�!�?W_�!O _�!-O�_�!UO�_�! }O�_�!�Oo�!�OGo �!�Ooo�!_�o�!E_ �o�!m_?/Q"q X/j  
OIASwb�� �������=� (�a�L���p������� ߏʏ��'��K�6� o���l�����ɟ��� ؟���#�G�2�k�V� ��z�����ׯ�ԯ� ��1��U�@�y�d���𯿚�ӿE*_DEV� K��M{C:۸̪f�OUT������?REC 1�,u��6� � 	� �Z�  
�j�m�w_Ìϝ���Q�bĽ��������w
 �Z�6 s��_�����@�Q��+vM���Y�鰕)�{�U*��B>����������ARߋ�+�,uж��r
ت���  UxR������z�K 鰝��a鰩���d�X���n�Ȋ�?nК��7�ߌU���R��R��R��E� �&� R鰟�a�=�[鰩���`�T���n�̊�*n�u����J�e��Hc�m��k� �  ���T���ե�z��.�Tp��n���6n�1zV�����~Kܽ�*i�(�t鰞�%���Q�QZ�� U�k���R�C���q;��~N@���e�a�*�P�Q>�Ɇ
D�鰱o��N���"��iR�b鰖R��RR������5/�|�� ��!UE���nм�$n�P�����*f�hR��Q��I͂*��J��_�沕C���nйB���/?/����I���P���f�./�Q<�Q�+�&$$�/,�/R/���&��`�m�R�W鰿T�/#���R�)[6?d��n����"^?�?������=�9 �?�?�?�?"OO2OXO :OhOjO|O�O�O�O�O �O_�O0__T_B_d_ f_x_�_�_�_�_�_o �_,ooPoboDo�oto �o�o�o�o�o�o�o :(^L�p�� ����� �6�$� Z�l�N���~�����؏ Ə����2� �B�h� V���z������ԟ�
���.��>�d�<�V� 1�I̜ �?����Eѡ�   -�~জ8��_T�YPE(��FZN_CFG �^������G_RP 2���/ ,BY�AY��_D;� Bq�A��B4�RB2�} �HELL�i������ ��<���%RSU1� Ͽ���>�)�b�M� ��qϪϕϧ�����߰��(�:�I��{ ���%I�w߉ߥry`%���%% ޤ7�_��d�ߏ�~�HKw 1Ō� �� =�8�J�\����� ����������"�4��]�X�j�|�x�OMM� ƌ���}�FTOV_EN��������HOW_REG�_UI��|�IMW�AIT��-0��O�UT��	TI�M��XVA�L-_UNIT�����MON_ALIAS ?e��? ( he��� �
.�6�[m �<����� �!/3/E/W/i//�/ �/�/�/�/�/�/?? /?�/@?e?w?�?�?F? �?�?�?�?O�?+O=O OOaOsOO�O�O�O�O �O�O__'_9_�O]_ o_�_�_�_P_�_�_�_ �_o�_5oGoYoko}o (o�o�o�o�o�o�o 1C�ogy�� �Z���	��� ?�Q�c�u���2����� ϏᏌ���)�;�M� ��q���������d�ݟ ���%�ПI�[�m� �*�����ǯٯ믖� �!�3�E�W��{��� ����ÿn������ /�ڿS�e�wω�4ϭ� �������Ϡ��+�=� O�a�߅ߗߩ߻��� x�����'���8�]� o���>�������� ���#�5�G�Y�k�� �������������� 1��Ugy���H����	���$SMON_DE�FPRO ����2� *SYST�EM*  �l��"RECALL� ?}2 ( ��}7copy �virt:\ou�tput\cal�prz.pc m�d: over �=>101449�728:9519O61  ��3���� }8r�tcp���</N/��:��_dv_xy.ls/�-/�/��/�Fr"� �'tp�v/�&�/�9?K?]?}	9r/�$z�/�,?�?�?�D�,z?�8�? �&9OKO]O��#!�?��+O�O�OaMtp�disc 0=>�laptop-3�jv248ms:?20980 �O�O�OG_Y_lBtpc?onn 0 �O_�_1_�_�_gG
xy?zrate �}_@�_�_�_DoVoiE!�W~�O13960 o &o^o�o�on@q�O�b�37224448�:878185 �o;M`NA�)!O�|v%r4��jD5�o _1,}�9�K�]���2	��-� ��Џ�O�O�n����;� M�`_r_��(���˟ ݟ�o/������<�N� a�s��~(���˯ݯ �� �����A�S�"fH6�� )����̿_��\test �/���=�O�b�#� �}z��/�����e���@�=����<�N�aM?r� Oz�ߣ�4�����j?�?�y��=�O�bLE �/�?~������oO��?��$s��<�N���C �?��M�߷������  �������GYl�~� ��+��as�� ��:L��� '���o���жG/Y/�";rfr�s:orderf�il.dat��tmpback\����c./�/�/d�2r�b:*.*�/�/�`�/��/H?Z?�w/ 3em�p0172.23�.254.7:17884 (?�?�?v�?}-r6*.d�? �=�?�?COUO�_4��?@O!O3O�O�Oi�ri�O �O�O�OF_X_k���$SNPX_A�SG 1�����}Q� �P 0 '%�R[1]@1.,7�Z?�h�%�_�_ �_�_�_�_.oo8odo Go�oko}o�o�o�o�o �o�oN1X� g������� �8��-�n�Q�x��� ��ȏ��������4� �X�;�M���q���ğ ���˟ݟ��(�T� 7�x�[�m�������� ǯ����>�!�H�t� W���{���ο��ؿ� �(���^�A�hϔ� wϸϛϭ�������$� �H�+�=�~�a߈ߴ� ���߻�������D� '�h�K�]������ ��������.��8�d� G���k�}��������� ����N1X� g������ �8-nQx� ������/4/ /X/;/M/�/q/�/�/ �/�/�/�/??(?T? 7?x?[?m?�?�?�?�? �?O�?�?>O!OHOtO�WDpTPARAM ��}U�Q W�	�xJP�D�@�hXOFT_KB_CFG  �C��U�DPIN_SI/M  }[�F_�'_9_�@pPRVQS�TP_DSB�N��Bu_�H�@SR ��[� &  AL_TC�E�_�D��FTOP_ON_ERR  �D��I�QPTN �U`A��RRING_PR�M�_ �@VDT_GRP 1ʝI�P  	�G�HZo lo~o�o�o�o�o�o�o �o# 2DVhz �������
� �.�@�R�d�v����� ����Џ����*� <�N�u�r��������� ̟ޟ���;�8�J� \�n���������ȯگ ����"�4�F�X�j� |�����ǿĿֿ��� ��0�B�T�fύϊ� �Ϯ����������� ,�S�P�b�t߆ߘߪ� ����������(�:� L�^�p������� ���� ��$�6�H�Z� l�~������������� �� 2Dkhz �������
�1.�CVPRG_�COUNT�F�8a�E\ENB'oW�M��D�_UPD� 1�[8  
E�B���%/ / 2/D/m/h/z/�/�/�/ �/�/�/�/
??E?@? R?d?�?�?�?�?�?�? �?�?OO*O<OeO`O rO�O�O�O�O�O�O�O __=_8_J_\_�_�_ �_�_�_�_�_�_oo "o4o]oXojo|o�o�o�o�o�o�oTYSDOEBUGf���`�d�pSP_PA�SSfB?,{L�OG ��ʱ�`�h  ����a
MC:�\XtYr_MPC ^}�����q
�� ��vSAV ��a}~t�r�e��wSV|TEM_TIME 1��W (B�>{�h�%�T1SVGU�NS�g'�����ASK_OPT�IONf������BCCFG ��G� @�*��`3�9A�j�U�g� ����ğ���ӟ��� 0�B�-�f�Q���u��� ��ү��ϯ��,���P�;�t�_������e ��ſ����
υ��@� +�d�Oψ�����}� ������������B� 0�R�T�fߜߊ��߮� ��������>�,�b� P��t������� ���հ�*�H�Z�l� ���~����������� ��2 VDzh ������� 
@.Pvd�� ������/</ */`/�x/�/�/�/�/ J/�/�/ ?&??J?\? n?<?�?�?�?�?�?�? �?�?�?4O"OXOFO|O jO�O�O�O�O�O�O�O __B_0_R_T_f_�_ �_�_v/�_�_oo,o �_Po>o`o�oto�o�o �o�o�o�o:( JL^����� � ���6�$�Z�H� ~�l���������Ə�� � ��_8�J�h�z��� 
��������ԟ
�� .���R�@�v�d����� �����������<� *�`�N�p��������� ޿̿����&�\� Jπ�6��Ϫ������� j���� �F�4�j�|� ��\߲ߠ��������� 
���T�B�x�f�� ������������� >�,�b�P�r�t����� ��������
(:L ��p^����� �� 6$ZH jl~����� � //0/V/D/z/h/ �/�/�/�/�/�/�/? 
?@?��X?j?�?�?�? *?�?�?�?O�?*OF�H@�$TBCSG_GRP 2�E��  ��HA 
 ?�  sO�OoO�O�O�O �O�O_�O'_9[LBSC��ZLd0 ��hQ?HA	 HBH�9XL�̈́V8TB   CyP�_�[xZ�_f�RD�_�]A��_pQ�UA�QTQ1o�Z�6ff�_^g@H@C��_�n@�^o�j	`C��o�o�o�n�_�oh Vh<uO,z��bt���{?Y����t�	V3�.00kB	lr;2c�s	**�"�pGB9��v�a�33H@\��y p�B�q��  ������LAJ�CFG �EedA g@����������� �5�C�@C�i�T��� x�����՟������� /��S�>�w�b����� ��ѯ�������=� (�a�L�^��������� ߿�kB�0��� �ʿ S�>�cω�tϭϘ��� ������+���O�:� s�^߃ߩ�HA4O��O ������(��L�:�p� ^����������� � �6�$�F�H�Z��� ~������������� 2 VDz��?� �`���
@ .dRt���| ���//</N/`/ r/,/�/�/�/�/�/�/ �/??8?&?\?J?�? n?�?�?�?�?�?�?�? "OO2O4OFO|OjO�O �O�O�O�O�O�O_� 6_H_Z__�_x_�_�_ �_�_�_o�_,o>oPo bo o�oto�o�o�o�o �o�o:(^L �p����� � �$��H�6�l�Z�|� ����Ə���؏��� � �2�h�V���z��� l_ڟ쟪���.�� R�@�v�d�������Я ������*��N�<� r�������b�̿��� ޿ �&��J�8�n�\� �πϢϤ϶������ ��4�"�X�F�hߎ�|� �ߠ���������
�� �T�Οl�~��:��� ����������>�,� b�t�����V������� ����(:��p ^�������  6$ZH~l ������� / /D/2/T/z/h/�/�/ �/�/�/�/��?"?�� �/d?R?�?v?�?�?�? �?�?OO*O�?�?`O NO�OrO�O�O�O�O�O _�O__&_\_J_�_ n_�_�_�_�_�_�_�_ "ooFo4ojoXozo|o �o�o�o�o�o�o0 @fT�?6?� �p���,��P� >�t�b�������Ώ�� ������L�^�p� ��<�����ʟ���ܟ �� ��H�6�l�Z��� ~�����į�د��� 2� �V�D�f�h�z��� ��Կ¿����.�� F�X�j�ϚψϾϬ� ��������<�N�`� r�0ߖ߄ߺߨ������  �� �����$TBJ�OP_GRP 2�����  ?��4�;���B����0�O���@�}� �� ���� ���S�	 �BL � ��Cр D�"�S�����?fff~��:lB ��߆ff@���33D  ���+��6�����h�z�����9�<�b�Y��?�٢������A�6��D��$�[��������
9�P�A���@����C��R�= ��UA6f�fhX�D/��z��͌�����a� 9�����@1��tz�&��{�3�33<T�8����?��?L� 9 S�B�Zcu�

�� >�ff�D���L^�^�%/ F8/"/0/^/�/j/$/ �/�/�/�/�/?�/�/�>?X?B?P?~?�?�C���1�5	V�3.00��lr2c��*�0����OG E����E�A E���E��3E�i�NE�!hE����Eۑ�E�I��E��E����E�rF��F�FM�(F�5F�BFaOF��\F"f$Bz � E�@ E��� E�� E� � E��@�� E}��@�� E�~@�Ԇ@�~@� F�   F� F�$ Fj` F��@ F�P F��` 9�IR9��o�<�ED:(��O
R�S��DI_0�ESTPA�RS�@��M�1�HR�cPABLE 1ْB�,P�NX#W (|�YNWNXNX�T�NW	NX
NXNXT�U�NXNXNX��A}SRDI�_L���_�_�_�_�_�U^dO foxk�o�o�o�o�n~R	SdoJ� (j��� ����	��-�?� Q�c�u���������Ϗ �'�cpg�\"� /A�_�_o#o5oGh�~R�NUM  V��L����� �@�@~R_CFGG �񛞓��@4��IMEBF_TT�iQ��J�vP3�VER��C4�I�3�R 1=�B�
 8O��ড ��-�   ������į֯���� �0�B�T�f�x����� ����ҿ����Q�,� >�T�b�t�s�_�`��@J�
4�MI_CWHAN?� J� �ßDBGLVI�A��J�3���ETHER_AD ?��3��K��τ�L�.���oROUT]�!B��!~Ԝ�o�SNM�ASK(�J�9�255.���3����0��OOLOFS_D�IiP���ORQCTRL �k��c_f�8U���� ����������,�>��}�z�L�^���_QPE?_DETAI�+��PON_SVOF�F!��P_MON� ��H�2��S�TRTCHK ��B�eߦ�VTCOMPAT��3Ӥ����FPROG �%B�%  AL_�TCP5���PL�AYjX��_INSWT_M�� �����US]�UgLC�K��QUICK�ME��!gSCR�E>+�tps�0g�Y^���o_s�PR	�SR_GRP 1�B�_ ؓ�.� ���/�3/!/W/E.�0�~/�*Q!��/ �/�/�%�??�/'?? K?9?o?]??�?�?�? �?�?�?O�?5O#OEO�kO	12345G678O�O^RXX�1��
 �}�ipnl/�@gen.htm�/�O_�_(_:_PpPa�nel setup>\}4~_�_�_�_�_�_ m_c_o"o 4oFoXojo�_�oo�o �o�o�o�o�o�oB Tfx��A7 ����,�>��b� ���������Ώ��W� i��(�:�L�^�p�� ����ʟܟ� �� ��6���Z�l�~��������+��UALRM�� G ?B�
  ͯ���J�=� n�a�������������߿��4��SEV7  ��f��ECFG �����ƍ!A��   Bȡ
 5ϡ+� ���������#�5�G�@Y�k�}ߋ�r�����C ��/��@�Ik?u�(%(��  �A�,�e�P��t�� ����������+����� ����9�I_�=HIST 1����  ( �c���%/SOF�TPART/GE�NLINK?cu�rrent=ed�itpage,,1 ����������
�(����menu��955����m�� 2D148?,2 _XY\�`���53��Z�w��*<��0f�//,/�'L�E34����4���/�/�/�,C/��CAL���/?"?4??/lQ/��71��MV�/�?�?�?�=�!��!� �?�?OO/OAO��? kO}O�O�O�O�OTO�O �O__1_C_�Og_y_ �_�_�_�_P_b_�_	o o-o?oQo�_uo�o�o �o�o�o^o�o) ;M�o�o���� ���?��%�7�I� [�m�p������Ǐُ �z��!�3�E�W�i� ��������ß՟��� ���/�A�S�e�w�� ������ѯ������ +�=�O�a�s������ ��Ϳ߿���'�9� K�]�oρϓϖ����� ������ߠ�5�G�Y� k�}ߏ�߳������� �����C�U�g�y� ���,���������	� ���?�Q�c�u����� ��:�������) ���_q���� ����%7� [m���DV ��/!/3/E/�i/ {/�/�/�/�/R/�/�/ ??/?A?�/�/w?�? �?�?�?�?`?�?OO�+O=OOO:
�$UI�_PANEDAT�A 1�����A  	��}  frh�/cgtp/wi�dedev.st�m[O�O�O�O�O�L)  ri�O&_A �@ >_P_b_t_�_�_�O�_ �_�_�_�_o(ooLo 3opo�oio�o�o�o�o��o :� � � p # Q�8_=Oas�� �o�._����'� 9��]�o�V���z��� ɏ���ԏ�#�
�G�@.�k�}�d���y�� �C�����)�;� ��_����������˯ ݯD�����7��[� m�T���x�����ٿ� ҿ���3�Eϸ�ʟ{� �ϟϱ�����(���l� �/�A�S�e�w߉��� �ߔ��߸������+� �O�a�H��l��� ����R�d��'�9�K� ]�o����������� ����#��G.k }d������ �1U<y�� �������	// n?/��c/u/�/�/�/ �/$/�/�/�/?�/;? M?4?q?X?�?|?�?�? �?�?�?O%O��[O mOO�O�O�OO�OL/ �O_!_3_E_W_i_�O �_t_�_�_�_�_�_o �_/oAo(oeoLo�o�o �o�o2ODO�o+ =O�os��O�� ����j'��K� ]�D���h�������ۏ �����5��Y��o�o}�j�����ǟٟ���)��"��u�N� `�r��������̯�� �ׯ�&��J�1�n� ��g�����ȿڿ������x�c�k�$UI_�PANELINK� 1��e�  �  ���}1234567890W�i�{� �ϟϱϹđrU����� ��)�;���_�q߃� �ߧ߹�Q�Q�
�����qS�  SOF�TPART/GE�N9�?CONFI�G=SINGLE�&PRIM=mainedit ���A�S�e�Q�
��M=�wintpe,1 8�����������.� @�R�d���������� ��������*<N `r
����� ���&8J\n �������~�� 0,  1� E5�or
�K.- co2/s/V'�/�/�/ �/�/�/�/�/?1?? U?g?J?�?���ߞ?�? �=R��OO/OAOSO eOX��?�O�O�O�O�O �OxO__1_C_U_g_ ���e�a�]�R�_�_ �_�_�_	oo��3oEo Woio{o�o�o.o�o�o �o�o�oASe w��*���� ��+��O�a�s��� ����8�͏ߏ��� '���K�]�o������� ��&'ӟ�t?	���� ?�"�c�u�X������� ϯ�����)�;��4 �]�_�?u_�?����п �����O*�<�N�`� rτ�ϨϺ������� �߃_�_�_\�n߀� �ߤ߶�=�������� "�4�F���j�|��� ����S�������0� B���f�x��������� ��a���,>P ��t�����] �(:L^͟ �������� /�6/H/+/l/~/a/ �/�/�/�/G��/k� ? ��D?V?h?z?�?�?�? ���?�?�?
OO.O�? ROdOvO�O�O�O�-� ?��__*_<_N_`_ ��_�_�_�_�_�_m_ oo&o8oJo\ono�_ �o�o�o�o�o�o{o "4FXj�o�� �������0� B�T�f�x�������� ҏ���e�,��/P� b�E���i��������� �՟���:�L�/�p� ���/��?ʯ9?� � �$�6�H�;Ol�~��� ����ƿؿg���� � 2�D�V��O�O�O�ϰ� ��������
ߙ�.�@� R�d�v߈�߬߾��� ������*�<�N�`� r���%�������� ����8�J�\�n��� ��!����������� "��FXj|�� ���e���0 TfI�m�� ����/��υ����s-�$UI_P�OSTYPE  ���� �	c"s/w/_QU�ICKMEN  ��+b/�/�!RESTORE 1���  ���"*?<?`9m [?�?�?�?�?�?o?�? OO&O8O�?\OnO�O �O�OO?�O�O�OGO_ "_4_F_X_�O|_�_�_ �_�_�_y_�_oo0o Bo�OOoaoso�_�o�o �o�o�o�o,>P b�����yo ���q#�L�^�p� ����7���ʏ܏� � ��$�6�H�Z�l��y� �����؟���� � ßD�V�h�z�����A��¯ԯ���
��'SC�RE� ?�-�u1sc%0uU2E�3E�4E�5E��6E�7E�8E��"UGSER'�,�>�T&��G�ksO���4��5*��6��7��8��� �NDO_CFG ��+  $0 �� PDATE ����Non�e V� SEUFRAME  $���$�RTOL_�ABRT/σ"F�E�NBP�A�GRP �1�9�!Cz  A��ä�	!�϶�����������?��� Up���_�MSKG  s�{�_�N,�%Y%|�%���߂"�VISCAND_wMAXq�I�[����FAIL_IM)Gq�^ �	 #{����IMREGNUMrq�
���SIZqӶ$0���,�O�NTMOUO�s�����N���d � ~����F�R:\�� � �MC:\P�\wLOG��B@�� !���������%�z MCV�����UD1(�E�X1�����TRAIN��^ o����)� (�!=��ͧ�������� ��������"4F�Xj|����PO�64_7����&3n6�I�LI��
��V���f@��� =	S�ZV���W�AI��STAT' ��	 @������$�/��H�2�DWP  ��P GC �"�2(9��A/��_JMPER�R 1�+
  ���2345678901�&���/�/�/ �/�/??8?+?\?O?��?s?�?�?�L�ML�OW����д�_T�IW��'��MPHASE  ����-@��SHIF�TM�1'��
 <�<��vOEUO{O�O �O�O�O�O�O _�O	_ /_h_?_Q_�_u_�_�_ �_�_�_o�_oRo)o�;o�o_o5E���	�VSFT1�uV��M�c �5���� �����A� W B8�`�`���psq�b�s]Ьg#ME> s����f	��&%�5AM������1��$�T?DINEND[�\؂�tOp�S߬wY��Sp��y�0q����G�#��F��&��x&���xRELEA�qϋtV�h�q_AC�TIVԉ|�
��A �ۗoV��
��RD� Տ�YBO�X �ｨ�������2X��190.0.�8�3����254��0A��� (�:�����rob�ot�d��   �pF�{���pcɐ����Ꝋ������a����ZABC
����,� %��⚯ O�5�r�Y�k�}���̿ ���׿�&��J�1�HCπ��Z9������