��   &��A��*SYST�EM*��V7.7�077 2/6�/2013 A�   ����DMR_GRP_�T  � �$MA��R_DO�NE  $O�T_MINUS �  	GPL�N8COUNP �T REF>wPO�OtlTpBC�KLSH_SIG�oSEACHMS9T>pSPC�
��MOVB RADAPT_INERP ��FRIC�
C�OL_P M�
G�RAV��� HI9S��DSP?��HIFT_ERR-O�  �NAp�MCHY SwAR�M_PARA#� d7ANGC zM2pCLDE��CALIB� D~B$GEAR�=2� RING��< �PLCL*w ��STA� >mTRQ_M���LINK"2&SX�<*Y<*Z/)II*IzW*Ie$ �RV*� L $� E�NBpV_DEBuU��!PNU;%�� UNEVEox��!8� �$�A�SS  �����!����� V?IRTUAL�/1�' 1 5�� ��� ��b?M?�?q?�?@�?�?�?�?O�>!L�M1HO6L�慄��}L�����b��KNY��_B5O�O1O[L��O�O�O�O�O_�K A_GR0_m__j_�_���d�_�_�_�_��=L3���_"o?�#o��@�Cohozo�o�o�o �o�o�o�o
.�_ 5YgwQ�4  2�_����� ��$�6�H�Z���< ���������̏ޏ�����&�8�J����$n% 15B1D�U5a�����_ ���_�ϟ��,�� )�b�M���q������� ݯ�����(��L�7� p�[�m�����ʿ��� տ߯!��H�߿l�W� ��{ϴϟϱ������ ��2��#�e�'ߌ�#� �ߛ��߿�������.� �R�=�v�]�gߩ�k� ��g�������<�'� 9�r�]����������� ������8#\G �k}����� ���1�X�|g �������/ 	/B/)/3u/7/�/3/ �/�/�/�/?�/?>?`)?b?M?�?[�RVk�r�`{?�?s?�?Hjx�?&O8OJO\OnO �O�O�O�O�O�O�O�O _"_4_F_X_j_|_�_ �_�_�_�_�?�_o�_ 0ooToOxo�o�o�o �o�o�o�o,> Pbt����� ����(�:�Ao^� I�n���{���ko܏�  ��$�6�H�Z�l�~� ������Ɵ؟����  �2�D�V�h�z����� ��¯�����߯�Ϗ @�R�d�v��������� п�����*�<�N� `�rτϖϨϺ����� ���	�&��J�1�Z� ��3��߶��������� �"�4�F�X�j�|�� ������������� 0�B�T�[ߕߊ�u��� ��������,> Pbt����� ��(:L^ p�������� �/�6/��Z/l/~/ �/�/�/�/�/�/�/?  ?2?D?V?h?z?�?�? �?�?�?�?�?
OO#/ @O+OdOvO]O�OM/�O �O�O�O__*_<_N_ `_r_�_�_�_�_�_�_ �_oo&o8oJo\ono �o�O�o�e