��  ë�A��*SYST�EM*��V7.7�077 2/6�/2013 A�Q  �����ABSPOS_G�RP_T   � $PARA�M  �  �ALRM_�RECOV1   $ALMO�ENB��]ON�iI M_IF1� D $ENA�BLE k LA�ST_^  d�U�K}MAX�� $LDEBU�G@  
GPCOUPLED1� $[PP_P�ROCES0 � �1��URE�Q1 � $�SOFT; T_I�D�TOTAL_�EQ� $,N�O/PS_SPI�_INDE��$�DX�SCREE�N_NAME {�SIGNj���&PK_F�I� 	$TH{KY�PANE7�  	$DUM�MY12� �3��4�GRG_S�TR1 � �$TIT�$I��1&�$�$T�$5&6&7&8&9'0''��%!'�%5'1?'1*I'1S'1]'2h"GSBN_CFG1 � 8 $CNV_JNT_* ��DATA_CM�NT�!$FLA�GSL*CHEC�K��AT_CE�LLSETUP � P� HOM�E_IO� %�:3MACROF2R�EPRO8�DRUeNCD�i2SMp5�H UTOBACK}U0 � �	�DEVIC#TI\h�$DFD��ST�0B 3$INTERVAL��DISP_UNI�T��0_DO�6E{RR�9FR_Fa��INGRES��!Y0Q_�3t4C�_WA�4�12HGX�_D�#	 d �$CARD_E�XIST�$FSSB_TYPi�� CHKBD_S�E�5AGN G�� $SLOT_�NUMZ�APRE�V��F�1_ED�IT1
 � *h1G=H0S?@f�%$EPY$�OPc �0LE�TE_OKzBUS��P_CRyA$��4�FAZ0LACI�wY1KR�@k �1C�OMMENy@$DGV]QP� ���+�BL*O�U�B , $��1V1AB0~ O�L�UR"2CAM_�;1 x�f$ATTR��@0�ANN�@�IMG?_HEIGHyAc�WIDTH�VT�CYU�0F_ASwPECyA$M@7EXP;$� Mf��CFcD X O$GR� � S!1zU`BfPNFLIC`<~d
UIREs3���AOMqWITC)H}cX`N.0S_d�S�G0 � 
$WARNM'@f�̍@� LI? �aNS=T� CORN��1�FLTR�eTRA�T@0T�`  $ACC�1"p '|�'rORIkP�C�k;RTq0_SF� �!�CHGI1 E[ Tz`u3IPpCTYVD�@*2 �P��`� 1zB*HD��SJ* ��q2�v3��v4�v5�v6�v7��v8�v9�vqO�$ <� so�o�h��s1�PO_MOR~. t 0�Ev�NG�8`TBA� 5c���A�����]@����ϋaP�0Ѕ*��h�`
P�@�2� �,p�J,p_Rrrqo@+�1J/r/�J�JVq@��Cj��m�g��ustP�_}0OF� 2  @� RO_���Wa�IT8C��NOM_�0�1ەq3���cD� �;����hP���mEXpG�0� �F�p%r
$TF�x�JF�D3ԐTO��3&@U=0�� e�H�24�T1��	E�� �e��f���f��0CPDBG�;a� k@$�PPqU�3�f):�L�A�AX 1�dUN�v$AI�3BUFuF8����! |�`��`PI��P�r�Mq�M~�䠁�F>r�SIMQS���G��QE�����MC�{� �$}1JB8�`S�}1DEC����r��:ܴz� ě0�CHNS_EMP��r$Gg�=Ǎ@_x��q3
p1_FP���TCh�@`�b��q0 �c}�y�G�� V�AԂ��!!���JR!0ԂSEGFRA.pv 7a}R�T_LIN�C��PVF������Y���Q��)B|����( '�� �f�e�S���Q��.0��p�B��A����SIZC�ћ�z�T��g���|���QRSINF3� �p����?�������؄����Lot��G�*�C3RC�eFCCC�`+� ��T�h��mh�SbA�� h�*�f��:�D�d�c2��C��PTA����0w@�撀��EV���jUF��_��F��N&��G�� X����r��1i��! ���,��hRGNP��0qF����R}�D���2}�LEWN��Hc6���C��K�uvqRcDx :�L��ou2���A�6N`Co�$LGp��B�1aP��s@�dBWaA?@���~0R����dME%`��d�f_RAs3dAZCh���z�OkqFC�RH`X`F�`��}��,�ADI;� 6b � ���`�p�`5cn�aS�@1�7a�AMP�Ē�PY8CU�MwpUt��iQU� $�P���C�CG1������?DBPXWO���=�p$SK��2�0� DBT TR%L�1 ��Q0Ti� �P�DJ�4LAY_CAL�1R !�'PL	3&@�0ED��Q5'��5'̡(�D�B��1!�W�PR� 
�1 0�1g" �PA$�q{$�� �L�)!#�/�#mp�0$�/�$�C�!%�/�$ENE�qr�&�/�#d R�Ep�"'H z�O)@"$LF3#$�#xB� W;���F�O[ _D0m�RO�(@���u��j���3R�IGGER�6PA�%S���ETURNܦ2RcMR_��TUr�`?�u0EWM���GN�P��zBL�A��E��$$P"#�CP� ��&@��"k�C5D�mpD�A#��p4\1i�FGO_A7WAY�2MO��fQ�g�CS_(<�QIS �����c�C���A�����B�t�Cn��A"�FW����DNTV@��BV kQ�����S˳W�sU��J&�U�� ��SAF�E�ZV_SV6bEOXCLUl�����'ONLA��SY��Q�tOTBa��HI_�V/M�PPLY_|�a��VRFY_#�q�Bd�_ )�0���_+�Ip � �TSG3� *�b݀�0 AA��a*����0��Vi.b%fANNUN� rLdKIDp�U�2~S@ �`mijarj�f�Rp�OGI�"+��$1FOb�׀OT@w1� $DUMMAY���d[!�d١�|& �E, ` 8�HExs��b�SB�$�SUFFIA�@ ��@�a5�g�6�b�MSW�E-{ 8��KEYI����TMZ1^ӌq�1�v�IN�����.{ D��HOST? !�r���t[ �t٠�tYp�pEM>���$�k��pL��UL���/ �|3��r��DT50�!0 � �$9��ESAMP��ԕF��������I��0��$SUB e�Q�� �C�:��G�SAV��r���G�C�� ˇ�PnfP$80E���YN_B�1� 0��DIad�@O����}$]�R_�I�� �ENC'2_ST � 2
ԇ J���L�q~S�`;�����!3�M�I��1|:�p�4  L�3�M��0�0K�4'a��AVER�q��}��M�DSP�v��PC��U���\ì�V7ALUŗHE� ���M�IP@���OP5P7  �THS ��D�6�S�F�F�³�dL�0�T��SC��Q�d:�ETo��5zrFULL_DUY�da�0��O�w��h�OT��A�0NO�AUTO�!6�p!$�\���cl�
��C�`�C����"��L�� 7/H *�L���n�b���$�0P�˴�� ֲ��[!���a��Yq��Tdq��7��8��9���0����1��1��1���1Ⱥ1պ1�1*�1��2
�2����U2��2��2Ⱥ2պU2�2�2��3
ʥ3��3����3��3�Ⱥ3պ3�3�3���4
�[���SE�"8 <��~��`��;I�����/��QFqE�0�0� 9 ,���Q? z@^ ?Q�А��ER@B#�8 ��@��� :�`�$TP�$V�ARI�<��UP�2�P; �pq�TD ��S|�1`3�����r�BAC�< T�pr��)��bP��@o�IFI)�@���$����P��rF�0��>� =t ;'�Ԡ��P'�ST(&�� @HR&�r0E����	%�C��	���_Cr�N��r��B��p�h�FOR�CEUP%bn�FL+US�`HN �E�h�RD_CMK@E8(����IN_��&v\Pg�REMM�F~Q���M �� 3
Kr	N0�EFF���N@IN�A��OV�Ml	OVAl	TR3OV���DT��mDTMX���m{@ �
��? �*[ ��CL��_:p']@$�2-	_
�;_T��X*
��@AQD� ��}��}!V1� �RQ��LIMIT�_�a椀�M��C9Lmd}�RIV	�a�n�EAR��IO*#PCC�����B�Bg�cCM@��R ��GCLF�G!DY�M(/�aR#5TWD�G��| s%�+��FSS& �s> �P�a�!r1��wP_(�!�(�!1��E�3�!�3�+5�&�GRA����?w��kPW晅ONT��EBU�G)S&2*�P{@a�_�E @�P�R� �TERMB5A<K5���ORIG0yBK5g@�SM_�P�r�G0CK5LED��TA�9DK6�PUP>B�E� -zAa��@.PY3.@A$S�EG�:f ELEUU�SE�@NFI,���2�1ޠp4�4B$sUF6P�$��FQ4@�wAG0T�Q�&�HSNST P�ATm�piBPTH	J�AߠE�p��2�P@؀	E)�؁��1R�@<�InaSHFT_��1|oA�H_SHOR �ܣ�6 �0$�7�@Dq�'�OVR#�na�@�I�@�U�b �QAGYLO=�z��I'"��oAj�!�j�ERV ��:Qh��J��OG @�B�0����U>���R!P"�ASYM.�"��1#WJG�уES�A�YvR�U�T @���E)�ᥳEP!�WP!�W�OR @MB��GR�SMT�F�GR��3laPA.@��`|�q�uG � ����TOC�1�`P<�@ �$OP���P�pՓá ��O�񖌀RE�`RC�AOX�pтpBe�`RmE� u�h�A��e$PW�R�IM�ekRR_p�c���qB H2�H���p_ADDR~��H_LENGqBPyqnq�q�R��S�I H��S���q0���u>Ӵu���u��SEȸ'�LrS��J� $��`��_OF�F��rPRM� ��aTTPu_�H�K (^p�OBJ?"ip��$���LE`C!�ȠL� � �׬�AB%_~TS�s�S{`��6*�LVN�KR��e�HIT��BG��LO�qt�fN�͂���`���`SS{ ��HQW��A�M�p`�INCPU�"VISIO�����+��t�,��t,��� �IO�LN��N̠�C^��$SLQb��oPUT_�$�`�{�P �V���F_�AS�"O��$L ��I����A��U�0�@�Af��`q�<PHY`���Ó�UO���#P `������ ڔ� �2�pP���`�(�L��Y�B��!UJ��Q�z�NEWJsOG-G��DISx�b[�K-�f�#R 
�rWAV�ǢCTR�C�ǢFLAG�"[�LG�dS ���Y�~3LG_SIZo����������FD)�I�4�E�*��D0 ���c$���𖶦����K���D0��� SC�H_��߅p�2��NT��F�T���E�"~�������U
�
�{`�L�	�DAU/�E�A�-��dE�;�GH��b<1��BOO��U�h Aɒ��ITp��y�[0ŖREC���SCR��ʑDI2ēS.@��RGO����˒����d�´���S�U���W�Ĳ�Ľ�J{GM$�MNCH,󾲑FNKEY%�KnM�PRGK�UFY��PY�FWDY�HL.��STPY�VY�@XY؀�Y�RS��H1`uۺ�CT���R��� �$�U	�m���
R��ݠғ`�G=��@PO�d�ڻŦ�M�FO{CUd�RGEX���TUIK�I{��� ��	������I�M��@A�S�`���@������ANA���2�V7AILl�CL!�U?DCS_HI+4`�D�s_�Oe�
!h�S���|�S����IGN 4��F�J��T�beç_BUj � V !PT�$*��rvD�Ϥ���a�!W �!Pi�'���0�1*?2?3?���_�>� X � i�=a0�5���Ņ�ID� tb	P5R�bOh ��\A�+ST	�RF�Y� �@~�  W$E�AC�y����8_�� Y L�؟0 ��@���`qFtǀ��FwҬ�_ Z �p����b���>0�C��[ �p CL�DP	��UTRQL�I{��T����FLAG�� 1�O�D������LD���ORG������hW>(�siT�r� 4\ ��#0��վ�Sy`T�0y ' �$�!�#RCLMC�$B/T/��)Q��!=1I�p_d]� d�RQ73$�DSTB�p�  � 6��-8AX�R |/8I<EXCES�b�s 5Mp�1^��D2�T 5��0_�p"6_A:&��;G?tY80K�d` \��GROU��t$M�B �LI9�CRE�QUIRDB�aLO�#KDEBUr�1L
YM��agb��`@�4C�"�1ND��`�c`b���̨�CDC���IN'��C��Z`���H��N��a#�� ��EPST�� �c\rLOC�RITp��P�Ap�1ޗ1ODAQ��d MX�ON�cF� R�fV�	X��b�U����w �FX0IG}G�� e �y @X�a��X�XR�Q%��Y	��X	��V<�0ғDATA$`�E�a��a�N��f t $MDEaI:�)Sf��^d�![g�H5P�@]ez��a_cANSW�a^d�a��^e�D�)ARz�� Xpg[ �0CU4�V�`��=URR2{�h �D2�`A��A�! ?d$CALI&0���GS�w2K�RINtb�t<�NTEg�(i�bCu��=RBqg�_N�qjPukr���$tht�2kuyDIV�&�DHi0jp+�l c$Vp�C�$M�$Z0R<!T 0R����b�emH ��$BELT˪ZA/CCEL���;�"�IRCO�݁m��yT���$PSi0
�L�ڰW��Cp�8��T�9�PATH���.���3]��Pl1�_<�r��Ł�"S C�r��_MG��$�DD�9���$FW�`7`���.����DE�PPABN�e�ROTSPEEՂ@L� JN�@���(0��$USE�_p�P&�ܦSYh>��p�! �QYN09A����OFFua��7MOU߁NGJ�܀sOL~�ٔINC�d�2Q��-2��� -2ENCSpa2U��,+4R�IN�I]�B����"n�VE��s^��23_UPօp�LOWL��[�` '���D>�2@Ep]�'��2C[pW�MOS����4MO��0�'P�ERCH  ��OV����蓼����� �$�8S+�� 2@����B��V�0^�O�L�0P��7O�U�UP"��������TRK��AYLOA�J��1���]�͵³3P� �RT1I�1	�� MO�O��-2�28 �`4�w�ٳ��?�pDUM2���S_BCKLSH_C]�P�ϐΦ� ���bn�"�y�Ñ���CLAL V��!���� ��CHK �SՐRTY����C�
�*!6a_�ä_UM�����C���SCL��W�LMT_J1_L< 0-օa:�E4�U�G�D�J�P�J�SPCd�ȑZ���3�PC �3�H_A@�2��C� cXT���CN_rN���.�S��%�V���:� ���]�9���C' �SH�r�*�*!9��9� p��^���9���P�A���_P��_ �"�Ŷ�!ճ����cJG����~�OG�׾,�TORQU��ON��޹*�B٢-�*�&L�_Wž�_�sj�P�sj��sj�Ir�I��%I�sFKP]�J�!��,c!�VC�0'42���1��{0��82��J�RK��+� DBOL_SM���"M�@�_DL�q�"GRV�q�j�sj�sKH_p��I���
COS��LN- ���� �p�	�p�	�����bFZ� ٦KMY��D�TH�eTH�ET0��NK23��s��s� CB�CB�sC&1n2�����s��SB�s��'GTS�1W�C.�2Q������$�'3$DU���8A!r��2P&�1Qb8V$NE�4�PI� ���"$%�v$�p�A��%p�'���LPH�5�"h��"S��3�3�3�"+3:2�pV��(V�(�p�,V�*V�;V;V";V0;V
>;VL9H�(�&�2�-�n�H;H;H";H�0;H>;HL9O�,OR�(O}I�.O�*O;UO;O";O0;O>;O2F�"�Y�T��'SPBALANgCE_T@SLE�H_�SPHq�hR��hR3PFULC�lX�R{W�R3Uz1i�
�UTO_����Tg1T2�Y�2N�� �`��Tq���Ps d���T�O�p!�L�INSEG���R�EVf��Q�DIF̨�zy1j_g�r1k�]�OBUa��t$yM�I`���SLCHW3AR>��AB��u?$MECH�TXˑ�a��AX˱Py�p�f�'�r�Pl 
�b�I��:�ROB�C�RW�-u�҈+��MSK_KP�tn WP �P_��R��r_tn���18�c�a�`_p`�y�_p�aIN:a��MTCOM_�C���po  �݀g`4�$NOR�ES��r��`�rp� 8U�GRJ��eS�D� ABג$XYZ_DA�!F�r�DEBU:a�q���p�q _P$��COD��� 1����`���$BUFIN�DXa�  !�M{ORRsr $�q�U&���u��ӑy��^��bGi�s � $SIMUL���8��>���F�OBJ�EjP��ADJUS<ψAY_I��8��D���s�Ԑ_FIב=s�TZ��c� ���`b�"�(�b`p0:G�D��FRIW�d�MTg�RO%�A�Eb����MF�OPW�O> Vpt0>�S�YSBU0[�$SCOP��I�����U���b`PRUN�rڕP�ArpDٖ�b��1�_�OUTΑ�a�t�$�IMAG��4\pv PDaIM��1��IN[ �0�RGO�VRDY�˒���P0�/�a�� L_�PB�}����RB�� 2��MkᜪEDb��` �N�@M��~Г��\�SLjPVpu x $OVSLfwSDI��DEX��@�q�����o��Vb��N�A��'��,��'�D�M~Ҥ_�SETK�Vpv @0U�^��ep�RI��j��
q�_�}�����q�^�dà*� w �H\q�`��ATUS><�$TRCx T��X�ѳBTMڷıI
��P�4}Ѱ���Vpx D\pE���β�0Ehbϱ�����ϱEXEհ����)�=���f�ym�]p԰UP��L�$�`6�XN�N���������� ��PG�uzWU�Bñ�e��ñ��JM/PWAI[�P��œLO7��pFA`���$RCVFAIL#_Cwq�p��R9��p��c��(�}�"�-�AR�_PL��DBTB8��,��pBWD ��p3UM*�"�IG�7��Qc�TNLW�"�}�Ry�iӻ�E�����|^���DEFSP` { L\p�`��q_��Ճ��UNI�����Ѐ�RD��Rb _ULA`Pͱ��P�pUq|-�#��q�O��tXPc�N�PKET��
��Pq�Uq} �h�ARSIZE�5p��=��u�S̀O�R��FORMAT��Pg�COנq�<bEeM�d����UX��<,�5p�PLIb�Uq�~  $�pP_SWI�`��/ G�~b�AL_ o�J��A�rB���C�r�D��$EL����C_lі� �� � ���r��J�30 �r��TIA4�Z�5Z�6�rMOM���f��s���pB��ADf��s����PU�NR����s���������Rt�� A$PI�&E�kq E�p-~-�-��WC�0$��&��9q�gE��eSPEEDL@G�����Ծ ����)�9����)�8�	)���SAMWPx�p0�1��MOVD� H$_S`Y%nk%_��	1�t�2�t����c��v��8�H�PxIN ����������(�+(+GAMM�<Vu!�$GETHE�U�ٓD5�
�POLIBRv���I�$HIu�_L�ݰpB�&E�(A�.� �&LW�-�&�,�)	6�&�1��f�`j��� ?$PDCK���"ٓ_�����E� ��b7��a4��a9�� $I��R��`D�c�b~�Ե`L�E�qkq���81��0�q6��`Vp�P/a?UR_SCR��A��r��S_SAVEc_D��8Ex�NO5�C��y�6�8@{$E�. {I��G	{I�@�J�KP �q��H� ���x" Mao���s���� d��6W2U�Cqy���:��M� �k�F� �aE��3�W<�@[�BjQWg@5r�U�R�R���Sc2jQM"��[C�L�W��M)ATr� ?� $PY����g$W`�fNG� O�`�b�b�b #�HЈ��a� ���c��%X�O���Z�e��ހRt� p䠰p�3+zO�O�O�O�O�a:5�_�r� |�E� 8@��>vs�>v��8@_�kwVvy�Eހu%�!sJB�\�P�"tP���PM&�QU5 �� 8*�QCO�U�1 �QTH#pH{OL<�QHYS��3ESe�qUE�p.B�Z�O��  q�P����%��UNְ�Q� ��OE��p� �P2�3��AÔ�R�OG�����Q2(�O�}�2������INFO�q� #�e���ڗRȾ�OI��� =(�0SLEQ�с �рi�C�{�D��L���`� OK0r���!E� NU!��A�UTTA�COPY�qu�?��`@ML�NHI�M�X�Cᐛ� Y�_RGADJ�q�i�X�Q��$ഖ�`
��W��P���0���l����EX8�YC0bI�ѪObp�q���n$�_NA9!��������`��� � Q���PORp�A�B�SRV0��)a�Y�DI��T_ ��{��������������5��6��7��8�y���S8BL��m�M�C_F�p��PL9A8An�ȰR��9��р���$iB����d� ,�0FL-`L�C@SYN�[�M��C?��PWRc��L���!�DELA��8Y�5�AD�a��Q�SKIP� ĴQ�4�OR`NT�� ��P_4��ַ@ lbYp���� ������Ƞ��ՠ���������9�1�J2�R� L�� 4*�EXs TQ%����(Q�����p�����p���R;DCf� �`��X9�R�p�����r���A$RGEAR_� IOT�2FLG0��vi��M%PC��B��UM_����J2T�H2N'�� 1������G8 T00 ������MlѺ`I��8�qREFr1εq� l�h��ENsAB{�(cTPE�0 �1���i�m���^Q B#��:��"������2�ҙ����������&�3�Қ7�I�[�Pm���&�4�қ��@���������&�5���1�C�U�g�y���&�6�ҝ����������&�7�Ҟ+=OPas�&�8�ҟ������&�SM+SK�q�|��a���E?A��REMO[TEF����a@0��(Q�IOQ5��Ic(P	��POW�0L�� �pZ�����#p%�L��U�"$�DSB_SIGN��1)Q%���Cl�(P%^��S232��b��iDEVICEU�S�,R'RPARI�T��D!OPBIT�`QY�OWCON�TR;�(Q��O'RC�U� MDSUXTA�SKT3N�p[0�$TwATU`PV"��0L����p_,PC�9�$FREEF�ROMSp��%�GsET�0�UPD(��A�2�PX P� J���� !)$U�SA^���6���E�RIO�P@bpRY$�5:"_>@ �P}1�!N�6WRKI[D����6��aFRIENyDmQ�P$UFw����0TOOLFM�Y�t$LENG�TH_VTl�FI1R�`-C�RSEN ;IOUFINR]���RGI�1ӐAIT�I��4GXӱCI�FG2�7G1��Ѐ3�BƱGPR� A�O_0~ +0!�1REЀ�E3�e�TC���Q�A�V �G8��"J���u1~! ��J�8�%���%m��5�0G4�OX _0)�L|�T�3H6��8���%r4JE3GU�W�P�W�R�TD����T��а���Q�Tm�$V C2����1���91�8��02�;2/k3�;3 �:iva�9=i�aa��^S�jR$V��SBVB�EV'�V�BK�����&c�p��F�"{X�@�2q�PS�E���$.rRC��o$AŠFwPR��Gv]U�cS'�� 7���E2I�G� 0�@qV`��p�d`���E0�@��=��
B5S!� �"�aRg����R�6�MN AX�!$�A�0�L(A���rTHIC´1Y���h�t1TF�EI��q�uIF_C	H�3�qI�G�a�pG1bxf���m���S@���_JF��PR��ֱ�S��Ԁ�Od �$SР�Z��GROU�̃TO�T�t̃DSP�JcOG���#��_P㱂�"O�����j��&KEP(�IR����@�M�R@�AP�Qn�Ep^�`�!�[�SYS6��"[�PGu�BRKP�B �.��pIq�p`��M���΂�`AD�!<̃9�BSOC׆��NӕDUMMY1�4�p@SV�PDE�_OP�#SFSP_D_OVR=���1C���OR�C�Nm0�F.����OV��SFR��pU���Fn��!#��C��A�"�LCH����РOV(�s0��W�@M��ĥF:�RO�#ߑ�_�p��� @@�u@VE�R�ps0OFSu@CV? �2WD6���2��ߑj2Y���TR�!|���E_FDOY��MB_CM�D�B�BL�b>�f��att�V"Q�240/p��N�Gg�z�AMx�Z�0���¿_M~��"7�����8$CA�7�D:����HBK81��IO�5���QPPA�=�"�M�5��͵���DVC_DBxC~� �3"�Т�!"��1��糖�3��� �pН�*��U�3��CAB��2VӆP�ѣIP��c�O��UX~�SUBCPU�r	�S�P P���90^S�Q׹c��."��$HW_C�Т��S��c�A�A�pl$UNI�T��l��ATTR�I"���	�CYCL���NECA��J�F�LTR_2_FI`_�G(��9&�1LP��?�>�_SCT�CF�_��F_��6��FqS8!����CHA�1��wᇲ�"v�RSD��4"����q�_T���PRO��>�� E%My_ܠ��8d��a� d��a��DI�b0!�RAILAC4��9RM��LOÐ C��Q*q��3q���+PR��SQ�pU��Cr�s 	�FUN9C��@rRIN'P�0�0��u��!RA��B� ����F�Ğ�W3AR~���BLQ�����A��������DA`����	����LD)0 ��Q1�q��*q1�TI2rQǁ�p$�xPRIA1�"AF
B�PP!|ߠ�<`8�R���MOI��A��DF_&@��51��L�M��FA�@HRD]Y�4ORG6 H����A�0 �MULS�E&@"�Q��a ��G�	�����$�d$�1$1� ���0���� xm�EG�̃�`cARހ��09�2�o��z�AXE�RKOB�W�A��_��œSY������SN�WRI�@s1���STR�� ��(�E�� 	%1��AB( �/&�a�ӰkOT0^�	$ߠARY�sf"���S@�	�FI��*�$�LINK���!��a_%#�%{q�"XYZ82�*�q�#'OFF���"�"�(%j B�j�4С��n�3FI��%7�q0���j���_J���8%��#�QOP_>$H+5�3�PTB\1�2�C��i�DU�&62�TURN��2r�5`t!}��p��|7FL�`@���m�0�%+*7�^	� 1�. K�	M�&82�Q�2rQ�#�ORQ��G��-( �+p��z�� 3q�E"��T�GOV�@-A��M*�y�4�E:�E@�FW�J��G���D�� o�*� ��A7�P�� y��E�A�GZU:ZU�C�G�ER���	6�E���B�TAFQ��)4�����r'�AX Уa2.q�c�W�c�W �c�W�p�Z�0�Z�0�Z %@�ZK@�Z��Z
!�V � �Y� 
i� i� *i � :i� Ji� Zi� ji�� zi�a�iDEBU{�$v�u��;q�0�"F7O�n�AB���6��CV�z� 
 fr����ukњw�!�w �!�w�1�w�1�w%A�w KA�w��\0��"3LAB"2|EwЄü҂�3 q EE�RVEN� �� $q�_NAǁ!_�PO����` �f�M�_MRA���/ d  T����ERR����~ TYi��RI�V"0�S��'TOQ�T)PL��T��ЅL�G�CJ /� p�PTl X���_V1�b�Q���
#�2�2+�����/@q��p��5�$W���V���VN�[�$��@�� �S���Q�	�EHELL_CF}GN� 5%��B_BAS��SR�vp0�K� �S���Jϐ1a�%Α2��3�4�5�6��7�8�RO0���� � NL:�3�ABn��АACK wv��)�o�u0i�n��_PU2�COq��OU��P��ӕ񰰒����TP�_�KAR�0��RE�m�� P����QU�E٩��@���CSTOPI_ALzs���� �TĠ�� S#EM[�w�k�Mw�y��TY��SO`��D�I���Є�=�װ_�TMK�MANRQ�ζ� E��$K�EYSWITCH���Ѱ��HE��B�EAT���EpLQE����&�U��Fd������SO_HOM�� O��REF�@PARi��R� ��C@�9O0�p ECO���>� _IOCM�4M��k������'�O�# D�!ۧH�U��;��M7��@�3FOR�Cߣ�� 􂰓O}Mq � @EtTxk�U#Po1B��O�o3B�4G�NP�X_AS��� 0�ݐADD��(�$�SIZߡ$VA�R�TIPr�q�G�A(ҷ��
�˨�r�t�n�SV�XC<����FRIF�R��aS%�7�x���NFѲ�EАO� x�PS�IڂTEC*�%CSKGL=�T�"�0&��V�D��>�STMTd
�o�P\�BW�@�?�SHOWw��P��SV� K�� ���A00�0�Q�� K���O���_���i���U5��6��7��8��9��A����6������20��F��
 �� ��U ����� ����0��� �J@��:�1G�1�T�1a�1n�1{�1���2��2��2��2���2��2�2�2� �2-�2:�2G�2�T�2a�2n�2{�2���3��3��3��3���3��3�3�3� �3-�3:�3G�3�T�3a�3n�3{�3���454��4��4���4��4�4�4� �4-�4:�4G�4�T�4a�4n�4{�4���555��5��5���5��5�5�5� �5-�5:�5G�5�T�5a�5n�5{�5���656��6��6���6��6�6�6� �6-�6:�6G�6�T�6a�6n�6{�6���757��7��7���7��7�7�7� �7-�7:�7G�7�T�7a�7n�7{�7ڈ�o�VP$�UP}D��  �Px���x�YSLO��� � ��հ�����QTAS�sTƠ���ALU}U����C�U��WFdQID_YLѳ�UHI�ZI�?$FILE_Σ�Tf�$u�_VSA��� h��+`E_B�LCK(�8bg�AhD_CPUQi��Qi����Sod_R1�ɢR ;��
PW,�d�[ �aLA�S��8�c�a�dRUN5��a �d�a�d��5��a�d�a��d �T�pACC����X -$&qLEN~�3t��&p䫠��Iѱ
�LOWo_AXI(�F1&q
�T2mwM��ɢ���I����Q�yTOR.�&p�{DW��s�LACE���&p�����_MAuйv�u�w�qTCV�|��wTڱ�;�1�<ѷt��H_��s��J����M��"ӠJ����u���u2q2��������s6�pJKцVK~��4���3ՃJ0����JJ�JJ��AAAL�����4�5Xr;�N1B�N���	��tL�p_k��#xo�"p��� `5`�GROU�PY�ӲB>$�NFLIC�ө�REQUIREv�EBUV�"q���кp2���#pɖ!qxг��� \��APP�RՐC���p
!�E�N�CLOz�,�SC_M ���A��u
!q޸�� 䣠MCp�r;�Xr|�_MG���C��,`��N��p��wBRK��NOL��t����Rϰ_LI��Hէ����JޠѤP� �p��p���p;��pD���p6�K��8��|������ Ғ�Mr:ql�Gqz�PATHv�������Rx��������pCNR�CaA��է���IN%r�UC�pwQ�Cd�U�M�Yop�����QE�:p�Gp�����PA�YLOAͧJ2L�HPR_ANqQ�L��`[�W�K�g���R_?F2LSHRё�LO\�䱕����ACRL_������޷C�XrH�P"�$yH���FLEX�� qJ%u� :2Dv�p4�K�GYq0�pPbt|F1Kљ� �׃�������E����/�A�S� e�w�����y���ф��@�蘏����J�ÊT���X����υ ��څ ��[����
�� �)���;�D�V�h�z�Y�J>��� � �������QIPAT��ё���EL4� �ؘJڿ��ߐJE��CTYRޱ��TN��F��ɗHAND_VB�p�ѹP`�� $�&�F2��K��ШRS�W��j��� $$M��}�R��E�� Uw�H��sA�PH����Q���A���P��A��Aɫ���j`��UD��DɫP��G�`�1)ST��9!��9!N̨DY�`���|� Y�鰋�KыǦ�J�ч�s�U�ХP��&��/�8�A�J�S�=��� ; �t�.R66N��/QASYM�����Ґ����Խ��ٿ_SH�����筈4 ��+�=�O�JV���h�'CI����_VI��dHN�u@V_UCNI�ÉD���J҅ �B�%�B�̦D�ųD�F �̓��������*Uc�I��-Y��H�`f��XQEN� �v�DIɠS�OwT8Y�YP��� ��I�1A��äQ�`Bc��S`�  p�a.a� �� ME�����R'R�1TkPPT@�0) ���Qz�~����0�Xa	iT@�� $DUMMY}1��$PS_�ЛRF��  ��Pf6�aLA��YP�jb��S$GLB_T >mU�e�PpQ p����Q� X	�ɗ`�SuT��ߐSBR���M21_V��8$_SV_ER��OÐL�c�cCL�`�bA5��O�RTPT O�P �� D �`OB���LO˰&uq9cp�`r�0�SYSq�ADR�TP�PTC}Hb � ,&����W_NA����tz�9SR���l =��M �u`�ys�u~�s� �s���������� �0�)�T�"�5�~� ��B����s�?�?�?D>Y�XSCRE)�p5�ȐST[�s#}�P!��t�Qr u_� Aq� T	� �`ob��a`�l��ҤԊ�g�c�O� ISb�c��UY�UE�TG� �ñjp^`Sq��RSM_iqmUU?NEXCEPlV֑XPS_�a����޳�p���޳R�COU�ҒS� 1�d�U�E�tҘR�b9�PR�OGM� FL�7$CU�`PO?Q��ִ�I_�PH�� �� 8џ�_HE�P�����PRY ?��`Ab_�?dGbOUS�� �� @�`v$BU�TT�RV`��CO�LUM��U3�SE�RVx��PANEԋ q��P@GE�U�<�F���q)$�HELPB�l2ETER��)_��m�A m���l���l�0l�0�l�0Q�INf��S�@N0�� ǧ1�����ޠ �)�L�Nkr� ��`T�_�B���$H�b T�EX�*��ja>�RELV��DIP>�P�j"�M�M3�?,iŠ0ðN�jae���U�SRVIEWq�S <�`�PU�P�NFI� ��FOC�UP��PRI8 �m@`(Q��TRIP>zqm�UNP�T�� f0��mUWA�RNlU��SRTO�L�u���3�O�3ORN3�RAU��6�TK�vw�VI�͑�U� $�V�PATH��V�CwACH�LOG����LIM�B���xv���HOST�r�!�R��R<�OB�OT�s��IM�� gdSX`} 2����a����a��VCPU_A�VAILeb��EX
��!W1N��=�>f10?e1?e1 n�S���; $BACKLAS��u�n���p��  fPC�3��@$TOOL�t$�n�_JMPd� yݽ��U$SS�C|6�QVSHIF ��S�P`V��tĐ�G�R+�P�OSURz�W�PRADI��P�_cb���|a�أQzr|�LU�A$�OUTPUT_BMc�J�IM���2��=@zr��TIL��SCOL��C����� ��Һ����������o�od5�?��ȦE2Ƣ+�0�T��vyDJU2��� �/WAITU����n����%��NE>u�Y�BO� ��� $UPvtfaSB��	TPE/�NEC ��� �ؐ�`0�R6�(�Q��� ش�S	BL�TM[��q��`9p���.p�OP��wMASf�_DO�rdATZpD�J�����Zp�DELAYng�JOذ��q�3 ����v0��vx��,d9pY_���9`7"\�x�цrP? ���ZABC�u� ��c"�ӛ�
  ��$$C�������!X`�P� � �VIRT���/� A�BSf�u�1 �%�� < �!�/�/? ?0?B?T?f?x?�?�? �?�?�?�?�?OO,O >OPObOtO�O�O�O�O �O�O�O__(_:_L_ ^_p_�_�_�_�_�_�_ �_ oo$o6oHoZolo ~o�o�o�o�o�o�o�o�{� ��AXLMT��s��#  ��tIN&8qtPR�EO��+vupXuL�ARMRECOV� �)XrzujF� �%�!d�������7�I�[�m�~��, 
�/��vNG�5� �+	 A�   ڏ�� PP7LIC5�?�%up�ՁHan�dlingToo�l -� 
V7.70P/36�v��
]�_SW2��D�F0j�W� 4�3Y�J�9�K�7D�A7?����
&�X��e	-�None���J����� ��T7�	���_��Viu�6s��U�TOz"�,tTy.�HGAPON� %��!z.�U��D 1�y� t�x�����y�.�K�Q 1�{ ) Hp������_ �����uq��"��" �!���Hեw��HTTHKY��"ٯ��� �u�����󿽿Ͽ� ����)�;�M�_�q� �ϕ��Ϲ�������� �%�7�I�[�m�ߑ� �ߵ����������!� 3�E�W�i�{����� ����������/�A� S�e�w����������� ����+=Oa s������� '9K]o� �������/ #/5/G/Y/k/}/�/�/ �/�/�/�/�/??1? C?U?g?y?�?�?�?�? �?�?�?	OO-O?OQO cOuO�O�O�O�O�O�O����TOĀ��DO_CLEAND�|��{SNM  ɋ���_�_�_�_o���_DSPDRYRL�_��HI!��]@�_ }o�o�o�o�o�o�o�o�1CU��MA�X �bTQNQS�sqX�bTB�o�B���PLU�GGb�cWo��PRUC4`B�P]klo�^�rO�r=o��SEGF;�K�+�6��_ �_}�������ŏ�0�LAPZom�/��+� =�O�a�s����������͟ߟ�6�TOTA�L�v�y6�USENUZ�g� HXL�NR���RG_STRI�NG 13�
��M,�S��
��_ITEM1��  n󝬯��Я �����*�<�N�`� r���������̿޿���I/O S�IGNAL���Tryout M�ode��Inp�B�Simulat{ed��OutT�OVERRW`� = 100��In cyclH����Prog A�bor^Õ�>�S�tatus��	H�eartbeat���MH Fauyl����Aler�� ���'�9�K�]�o�8�ߓߥ� ^S�� ^Q��������,�>� P�b�t�������������(�:���WOR9���r���L��� ����������* <N`r����8���PO���� ���9K]o� �������/ #/5/G/Y/k/}/�/DEV� -�/�/ �/??)?;?M?_?q? �?�?�?�?�?�?�?O�O%O7OPALT ��^A��8O�O�O�O�O �O�O�O__(_:_L_ ^_p_�_�_�_�_�_LOGRIxp��avO�_ *o<oNo`oro�o�o�o �o�o�o�o&8 J\n�_*�R�ݦq o������(� :�L�^�p����������ʏ܏� ���PREGbNK��$�r��� ������̟ޟ��� &�8�J�\�n������������$ARG_�r�D ?	������� � 	$�	+[�]���.���SBN_CON?FIG ��L��K�F�CII_SAVE  ��k�b��TCEL�LSETUP ���%  OME�_IO��%M�OV_H��¿ȿR�EP�|��UTOoBACK��V��FRA:\�8� �8���'�`��8�c�,�INUIa@8�^�,�?MESSAGz���������ODE_D��}�C���O� ��,�oPAUS!���? ((O��J� \�F�|�jߠߎ��߲� ��������B�0�f��t�%�*TSK  �5ݒϕ�/�UPD�T����d����X�SCRDCFG �1��� �������&�8�J�\� n���\�n�������� ��"��F��j| ����/e�2�GROUN����_UP_NAܰ��s	2��_ED���1
��
 �%�-BCKEDT-`��}��p��Pg3�p8�/�/�8���g2���E/��/��/~/��ED3n/&/�/J/�\.�/"?�/�/ED4 ?�/?�/\.[?�?5?G?ED5�?n?#O�?�\.�?jO�?�?ED6 ZOO�O6O\.�O_}O�OED7�O�Ok_�O�\.G_�_!_3_ED8�_�o�]-�_Vo�_�_ED9Fo�_�o�"o]-�o�oio{oCRoY_Vh�]1��{� LNO_D�ELGE_U�NUSE	LA�L_OUT �V��WD_AB�OR���~�5�IT_R_RTN�ǀH�ONONS)Ю������CAM_PAR�AM 1����
� 8
SONY� XC-56 2�34567890�Y �f�@����?�W�( С���8�h�х�ڎ��HR5ǃ��	���R570�B�Affފ������ڟ� ǟ�"���F�X�3�|����i���į!�CE__RIA_I����5��F��;�Я� ���GP 1]����s�����V�C󠸾�����CO�C ��(���ǀC8��@��H̺�CCX����Ch꺰p��x���� +C�����Ⱥ���+�=�G��ށ��HE>/pONFIG=�f��G_PRI 1�B�$r�����������(�~�CHKoPAUS�� 1���� ,wuj�|ߎ� �߲����������� 0�B�T�f�x����D�O���T���_MORGRP �2?� �\�� 	 �,��P�>� t�b���5�����eҒ.�?a�a�����K(���d�P�V��a�-`�/A�

s��������b&�i��ܦP�DB�����)
�mc:cpmid�bg��:� � +���p��U   �*�m�n3� ���d�~��~���{C�e��
�{g�+/�n��~f/s/i�u/�
?DEF �(K��)�b buf.�txt�/�/��_�MC�����d(,53����ʇ��Cz  B�p�B��Z�B�X�B���~B���B�<�C3��
�q�Dv��D:��"Df��DRt��DStD�a���=F�pgF=�C�Fi�WF��EF�2?Fj�I�	ބ	6��N��4���(D)~�2�/��ʄ3@9à1/  TB�{D�V@a  EI��5� F*� �F�G$ˀF[ߺ GR�kNGl���G��G���&H��G֟��H��߃]���  >�33 ��ށ�x�@F߂5Y�Ed��A���=L��<#�
 ��_�*2�RSMOFS�ظ.^�9T1��DE' ��L#
 Q�;;�P  0_*_^>TEST�"__���R���#o^6C"@A�KY��Qo2$I��B�0�� �C�qeT�pFPROG %�S�o��gI�qRu����dK�EY_TBL  �6��y� �	
��� !"#�$%&'()*+�,-./01��:�;<=>?@AB�C� GHIJKL�MNOPQRST�UVWXYZ[\�]^_`abcd�efghijkl�mnopqrst�uvwxyz{|�}~����������������������������������������������������������������������������q���͓���������������������������������耇��������������������E��`LCK�l���`�`�STAT�c_A�UTO_DO���O�INDT_ENB;���R�QY�K�sT2����STO��~��TRL�`LE�TE�ފ_SCREEN j�kcsc 	��UπMMENU� 1i  <�l�ol�K�u� ��FS����柽�ϟ� ��R�)�;�a���q� ��Я�����ݯ�� N�%�7���[�m����� ��ɿ�ٿ�8��!� n�E�W�}϶ύϟ��� ����"����1�j�A� Sߠ�w߉��߭߿��� ����T�+�=��a� s����������� >��'�M���]�o��� ����������:�#p)+�_MAN�UALӏ��DBC�Ou�RIG�$�DBNUMLIM��,1e
�PXW�ORK 1k �_-<_N`r�wTB_�  m���Y0�_AWA�Y��1G�@b=�P�_AL� =��B�YҀ��`�_� � 1!�[ , 

:&d2/o/�&J�Mt�IZP�@P��#ONTIM�M�d��&�
�e�#MOTNEND��o$RECORD 1'kU2)?�!�O�?1-?&k�k? }?�?�?88�?�???�? c?O*O<O�?�?rO�? �OO�O�O�O�O�O_ �O8_�O\_n_�_�__ �_%_�_I_�_o"o4o �_Xo�_|o�_�o�o�o �oEo�oio�oBT fx�o��/� ����>�)�7�t� � pu�����-��͏ ۏ�����N�`�Ϗ�� o����)�;����� �8���\�˟ݟ���� ;�Q�گI���m��4��F�X��TOLEoRENC�B�	"��L�Ͱ CS_?CFG ( +x'dMC:\���L%04d.CS�VY� cֿx#A V��CH�z _/�x.�G��},��RC_OUT )��- z/��SGN �*��"��#��08-JUN�-25 13:5�2��27-�MAY��4:38��]� Z�t������x.����pa��m��PJP���k�VERSI�ON ��V2.0.11~+�EFLOGIC {1+� 	d���ٓ��p�PR?OG_ENB�2���ULS�' ��p�_WRSTJN� ��"�EMO_�OPT_SL ?�	�]�
 	�R575x#?�74jD�6E�7E�50i�d�o�2E�d��j�"�TO  .����k�V_� EX�d��% �PATH ;A��A\��M�\_�~+ICT�F��, '�`��eg��}�STBF_TTS�(�	���Eм`���� MAqU��ߧ"MSW���- )��},t���.�!��]l�R�v������4SB�L_FAULy�/���#GPMSK��ߧ"TDIA��0؍���`���!�12345678#90xS�l�P�� ���//%/7/I/ [/m//�/�/�/�/�/�L0PV � ��/�2?X?j? |?�?�?�?�?�?�?�? OO0OBOTOfO8<x�gUMP$�I� ��ATR>�O�@P�ME���OY_TE{MP��È�3��84��DUNI	�w��YN_BRK �1��x�EMGDI_STA	��_�LP�NC2_SCR 27[��_�_�_ �_�&�_�_o o2or�nSUQ13y_+?|o�o��o�olRTd47[�Q��o�o���_> Pbt����� ����(�:�L�^� p������� ?Ǐُ� 0�,p��+�=�O�a� s���������͟ߟ� ��'�9�K�]�o��� ������ɯ����� #�5�G�Y�k�}����� ��ſ׿�����1� C�U�g�yϋϝ�ׯ�� ������	��-�?�Q� c�u߇ߙ߽߫����� ����)�;�M�_�q� ��ϧ��������� �%�7�I�[�m���� ������������! 3EW��{��� ����/A Sew����� ��//+/=/wa/ s/�/�/�/�/�/�/�/ ??'?9?K?]?o?�? �?�?�?�?�?�?�?O K/5OGOYOkO}O�O�O �O�O�O�O�O__1_ C_U_g_y_�_�_�_�g�ETMODE 1�5'Efa �t|�_GgRRO�R_PROG �%�Z%���HogTABLE  �[�1O�o�o�o�ZRR�SEV_NUM ��R  ���Q�`a_AUTO_ENB  u��SZd_NO�a �6�[�Q�b  �*�6p�6p�6p�6p�`+5pOast�HIS�cXa�P{_�ALM 17�[� ���6|6`+ t���&�8�J�x�_�bp  �[�4q�R���PTCP_�VER !�Z!�6oZ�$EXTLO�G_REQ�v�y�SIZ�܄T�OL  XaDzޘr�A ܄_B�WDo�%��fQ���_�DI?� 8'E�t�TXa b[�ST�EPg�y��P��OP�_DO�v$v`F�EATURE �9'EQ��Q�Handling�Tool � D�ER Eng�lish Dictionary��7 (RAA� Vis"� Ma�ster���
�TE0�nalog� I/O��p1�
0�uto S�oftware �Updateb� �"/�k�matic Backup
��d
!��g�round Ed�itB�  25L�Camer�aT�FX� "Loμ�ellT��L,� P��omm9�syhۡ�h600��scou���uct���p�pane� D�IF���tyle selectѡ;- /�Con��9�?onitor���Hd�tr�Rel�iabT�ϣ(R-�Diagno�s��Q�	�H�Dua�l Check �Safety U�IFc�Enhan�ced Rob �Serv��q ��v	ԸUser� Fr���T_i��xt. DIO� f�fi�� )�\��endܰErrzu�L��  prנ�*�rO�� @���E�NFCTN /Menuİv�����.fd`�TP I�n?�faco�  �
E�G��p;�k Excذg�C���High-Spe�ܰSki��  P�ar+�H���mm�unic��onsn��\ap��urf��?�X�t\h8�U���connZ�2�Т !�Incr���str)�8��M�-6�KAREL Cmd. L���ua��}��B�Ru�n-Ti�EnvB�(<�@�I�<�+��]s��S/W�"H��Licens�e���� ad���o�gBook(Sy�>�m)	���"MACROs,�¿/Offse\�fĜ���H�!�Y�M1��MechSto?p ProtZ�3�o 5
�Mi4��Shif\��B6S�MixܰQ�����H�Mode S�witchY�MoTk���.�� ��Mt�Q�g�� �5��ulti-T�������)�Posj�Regyi>���  ! �}PA�t Fun1מ�6iB/��R�NCum�Y�3�G�P/�|�� Adju���	�/2HS�)� yo(�8�tatu����AD ��RDM�ޱot�scove&� #e�v�㱗���uest 86�7.��o�\���SNPX b��Y��Þ)�Libr%�
�r't I���� "���Ҫ�.S�o� ��s in VCCM����� j������㣀/I�� 71�0�TMILIB�X����g�Accܨ���C/2�TP�TX�� �Teln���Y@����K�PC�Unexce{ptܰmotn��� ������\m725����w�5����  h640S?P CSXC�i �� j*�� RIN��We���50,���vrl�زme�n" ��fiP-�a����P��Grid�{�play F �O/��? ��ELR�;�|�20��OR�DK�sciiw�l�oad�41d�s�t�Patd��C�ycT�h���ori�ɰ:�7c Data&� qu6�2�0�*�p������FRL�amc�K�HMI �De��(����k�P�C�φ�Passwword�644���Sp�����D#YELLOW BO�	�?1�Arc%�vi�su����#ti�OpX�^�! 2��aO��po�� t��ֶT11o�����HT���xy�	�   $�t۠ig��10�Ơ 41\+�JP�N ARCPSU� PR+�8b!O�L0Sup�2fi�l� �!��E@-�;�croc�82��v���n$ 12jSS0]e4�tex-� I��7�So��tf�ss�ag�� e��У�P���,��� "Tc VGirt��v�!�����dpn�
�J3ނSHADf0MO�VE T�MOS� O TԠg�et_var fails l�>PU�~1E���� Hol�d Bus %�h���VIS UPD�ATE IRTO?RCHMA A�{��vYWELDTV S� ]�DtS: R7[41��ouiPb}��y��BACKGR�OUND EDI�T "RC$REPT�CD CAN C�RASH FRV�R 62z1�SCr}a��s 2-D���r ) "��$F�NO NOT R�E��RED �` �m ��JO� Q�UICKaPOP �FLEN m41�S�Loc��gRTI�MQ%�#�FPLNs: FG��pl m��r`�MD DEV�ICE ASSE�RT WIT P�CV;PB�AN#aA�CCESS M �.pc��Jo��Q�ui±�Kbldm�gUSB$ ��t & remov��� Pg�SMB N�UL� ;a|�FIX���C��ACHIN�,QOL�`MO O�PT ՠa��PP�OST0�WDU �C�wQAdd�`aYd���0io�2��k$P�`W\0.$0`�O�IN&�P:f�ix CPMO-�046 issu5eC�J/aO-�0�r7130Т- ��vR�SET VARIABLES-P{��R�3D m��vie�w d��M��&�e�a���b��of �FD�5P:N@x �OS-1y0`�h isc���t��s t�3lo��7 WA�PZ��3 CNT0 T��/"�ImR�)�c�a �Pu��POT�:Whenapew�B�STY E�{1t���ptKQdo G�ET_�p �p��V�MGR LOl�REAd0C~QW�~1��(�l�s�gD�ECT�pLpING IMPR�DR(p+PB�PROGRAM�E�RIPE:STA�RTU� AIN-�;�ӠM/ASCIyIzPÂOF Lq��DPTTB: Nv�pML$me P����`:x�mo&�a�llW`!�ӤTorBc�A�U�HC�iLp�Ըth�`n�@ c�h��/GEA�!�toyu͐�RCal���k�Sign`� N�D�ԗThresh�123��`��09p : MSG_P��+0er  �Q�Aܠzeron��0� H85��RImlA�n�2D��rc�0�I��OMEa`�pO�NaP5�  נSRGEG:FF-Д� ]�|'���KANJI���n��J��c�0asn� d�!OA imm�c �INISITALIZATI�����~1wem����d}r+� LB A�U�Wqminim�r�ec[�c!�R���m>$�ro -1>ѮS�ܰir��@ұJ�1pdETw�� 5`?�I��ow u��< se� 1lc��YbPM ���p�Q���R`vR&��lu\�3�Re 0��4q�q1#���m <a�arn��ঁ?Box fo��*PORWRI�PW�S���v�09 F�pup~�de-rel2 �d�p� j��`━b�etwe��IND� Q���igE s�nap|�us��s�po TME��T�PD#�DO�p#aH�ANDL 1\kP�`vR��ȀD�ny��S�v�Yopera�bil� �T*�: IH � l\p��Vq�Hb�R�< p�a*�c&2�O�`FA,�.�-QV�7. f.v��G-T�pi�s��� �ɠtmLine-Remark ^�� RM-�` W��#SPATH SA�+PLOOS UIqFc�+5f fig�pGGLA����Vrp�������U�0ther|�V� Trac��"�tW�\b�s7��d��t�� n�@  ����3:���dK�y���it k8�d�P;ayR![2]�ü�1: g��s��d�ow�XQ��0IS��q�qEMCHK ?EXCE C���OMF +�Xah�� 35\k��)���QBt���'b���2[�c���e �`k�<�S�� BUGr�:�cD$`PETp����f�c4��0XPAwNSI��DIG���@OoPmetTCC�RG EN��CEOMENT�A M̀�K {�`H GU�NCHG �`� ECXT�P�2�bQS��93 wP8�x�OR�YLEAKq  �H5gyq�PLC �WRDN R �O9 /u�QSPE=p��G*�V ��$�t�n720\3pGRI��A�rT�PMC� ETH��pSU<7p�`  j5/n�/PENS�PN,���*P ont�`BR�OW�`!sRMV 7ADDz CN q�DC���PT3 A�LA2@ ���pSV�GN EARLY8�R��ŰH57�Ga�JLAYҀE 5(@M�PPD�p*@�H�S I`P�OGUCH8���V�F�q��comH�x ��E�RROR� DE �nJ��RO�CUSRS8pI��N4<q�-158n7�ORSR xP#aUp�P��Rqy�T�Fz��;�pk��t�� g�Ղ�B�SY RwUNN�  a�`��BRKCT�!RyO�p3@ \apS�Ƣ�AXxP���h8x+ q��ISSUrp} sPX�PTSI��K1M10_�IP�SAFETY Ck�ECK[��Á�������<#X�� �T�WD2�@�@�IN=V��D ZOp�5�X��t�DUALy� "M6�0�"r�F#�E��dPdNDEX F�t*UF�"Pʀ�0s�FRVO117 �A�PT6�KtqFA}LPTP2477D�6_�P�!;HIG�� CC�t;SNPX� MM��tq�d~�Vq�q#�
"��DETEC�Tq*@RRU�qA�P�5p
�9 y�)<9���7�T��Pds� �k�	���!Q����� t\4A�;A0�27 "Ke@" 8@HI��qXF8@4@H�PRDC"�
�aMB8@�IXF�b���zOX@8@����a�G}E�B�Ccsc�r�J8@�Ndctrld.�A�NZE�A5�I�Q��!�`�Df8@\�`m�878�Q-;� ��� rm`�
���PR̠78�@RaI8@0q�Q (~\�Mp��0t��!{B8@\PtQ<OX�St0�3hB�3nO�Vtp�A�@L�CF�L��� �Rplcf���J8@�WTa�mai�E8@mubov2_miTA�O�S8@U`�T[tT�AqPr674�xSShape G�en��8@j�I�[R��`�@8@T����%q 1(u8@��II�^�Q�~C�a�[8@;Ynrsg:0�4� � 4�CtMSr68@�r5hB5�z�Vnretsp "�r�Po�wng0bGCRE�Ka�ޠ��DAT�E�k�cr�eat.�q�M�a��oksqgtpadx1P��(�tputZj@�{�������܆28@`����Q����sl�ov��� �hexH��TB�8�ď�keyH�8@�pmZb�NR�1u7A+�nrgc8@UQ��pp�bUZ�dp0aj�921xSpl.Collأcq�\A��R1Nq�UA� (J�8@ip�_�WA��_�Y���a7hB7�ͦtp~[� "TCLS9o<Kb��clskyh[:��s�pkckZd� ��$�TQ���dA�rx��710a- KAR�EL Use S=p�FCTN9�a�a7l�0s0a�� (�� �a��~C8@��MI��c�8hB8"   ��8@ v	��v	   lomatea99�q�M����E�mcclm5�CLM;�� �j̕�E�et���aLM�	�h�yasp,���mc_mot�B�N��`8@H����Q��su'���Q�ȕ�䅮���jo�i#�ߕ��A_loqg�Z���trc�B����ve�ϓ�v��Q�WX��6�finde�rxSCenter� F1�lSw520���ha6rX� (<�r1,�Q�Ձfi�Q � NH0�I�ۡ���A8@uL���tq�a "FN�DRVϳ���etgwuid�UID�C 8@���������TA@�nuf;��P���ƞC�B��_z�Ӡo��q�G������l���fn�drTY��2䁴tcyp"�,qCP MF�:}38@517��6s38�E��gf6�� (��K��Q��-�X��A&�tm6�P�İ ��Q���	�͘���tm�Ĵ�b8@e0j��TAiex��aP��Aa�ذ�cprm�A��l�_vars��
��dwc7 TS0��/�6��ma7AF��Group| sk� Exchang�J 8@�VMASK �H5�0H593 MH0aH5@� 6� +58�!9�!8\�!%4�!2���"(�/�@�;OMI� `@a0hB�0�ՁU4U1#SK (x2�Q�0I�h��)��mq�bWzR�DisplayImQ@QvJ40�Q8aJ�!(P��;� 0a��0�Ϙ� 40;�qvl "DQVL�D쌞�qvBXa`�uGHq��OsC��avrdq8�O�xEsim�K40FsJst]��uDdX@TRgOyB�Bv40)�wA�~���E�Easy �Normal U?til(in�K�11 J553m��0b2v�Q(lV40xU)���������k98�6#8Uϕ�|�rP "NOR��dw d.a}oKksu�O�W���O�Y�W`�j0�6�H� mOenuuyP6�M�`�wRX�R577V�9{0 �RJ989}��49b\�`(�fity�����e�<?L��Vsmh`��8�� C0�Sv�q�8����w�pn "MHMN<��ޣx�Ay`�o�3@�u�`f�І�x�t���tRzQ��LV��vP�tm���|I�1{oPx ��2|���I�3I/B�ogdstǏًmn吼���}ensu_�L<���h!!��Rt��?huserp��0���ʐcM�_l�xP�oxe��рpoper��|��xdetbo/� l>�x���Ps$p�`����OPydspweAb͓��z'R��u�Rr101&S՟{t�`12�Z4�30���D���`4�
�4�5���KQ�m[T��dUCal G40`�Q)p40}������9;��DA��� v	LATAu�mpd�\bbk9�68��68c�fb\l�41969y�9�|��D���bd� "B�BOXêM��sc�hed����m�se�tuM:�����ff ���40��n�41�ϒ�40q�col��|�1�cxc�ؘ���li�� X�0���j��&�8�4 �<�ro5�TP E��#��ryK42�r��;�(T+Q �Rec'�ʈ1Iw�84������Ak971���71�;���parecjo��QNS��[T���dXrai=l| nagek�M �,QT2 *� (�ĜR%<x�80!�bh��p��4��4��yDgl�paxrm?r "XRM�g�l�brf{���n����kl��9turbs�p��㧑- �l0195	�g�625C�M h�+���)89��	+��B6��o�ҹ���x�7�q40����pd "TSPD�=<��tsgl��l��:dQ���8Bct���K�vrE�aܮ�����  c�!���21�`�( AAVM l�2�0 �@fd �TUP him �(J545 �l)�`8 616 �%�VCAM ���CLIO �(�0:�5&  {(F\ MSC �R�t"PBsSTY9L�D!28 :2\ �NRE F2h SC�H6pDCS�U tpsh ?ORSR �rD!�04�SEIO�C& \fxh 54�2 LEX"� E�SETn�8!H ��s�h8 7H �M'ASK�Ø"7>���OCO*`x�!03P"6�!/400:66$ �G639.6[8LCH�!6OPLGR703�
5MHCR��0CЄ (! �06�A.f�8!54
��00DSWb 588�180 ��h!37 88 (%D�"02C24���2'7 q9�25��2�-6�05��9P�RST bBFRDMES�!zB��930 _ NB�A  6� HLBo 3 (~!SM�@� Con� SPV3C �8!20z���TCP aram�\TMIL �A��@PACETP�TX �@p TE�LN 96��29^�%UECK��r UFRM et��P!OR ORP IP�L%CSXC�0j��1CVVF l �FQHTTP satA")�I#� CGHP�8ZIGUI��0�hPPGS T�ool� H8�@d�jZ��!@�h!63��%�@32Q\�31 �B�h!96�%R65�1�Rs�!53 T7FAD�R41�8"[1 ��oo�"9��41775�"/@�P�VCTO�@�U�!s�h!80�%PRXY<�R�!770 �b8 ?885 ol3P� L� аdi� �`ڳ�h LCP{Q� TSS �b�26:����@�CPE �HT@V�RC~�tQNL <��@002 %��b�	0dis� �`7 `<��a\0�T�`1 �`{en�b4 652�`)FU02Q0Πo`dp�Ptu�r4 $�r5N��RU0p@n�se�QJp1 AP�FI[ Jp3�g34>�g40 alxrlE1t44w46� ts U0  7v�0�O��r5�e�p7 po "sw�a61:���r4��r5 QpwGr`�$�p8R�"sP`�tQ�b�36w77��w8`�v83���r8��&:��pOq8�8 "/rkey8�9F��a;90�91 p�#@���� �D095�g9-7*pur�A1@d����P|P�q1�0Qpl�Sq1p#4��]a!s1&@sl༂8�Ӽ�$\1�d1�`��v�@�{�14p�ae��5 �h2��`�6ޣ��7�f1p@��d�YpCqd�ـd�1�`uq��� BCu1< Oq� ��7ReU1$ �u1�Pϱ� ܺ�@- WQ158 ase C���9 B��60 8�2ń�p���4 (Wai��`吢!��i7E��8�EU1P`�ro9�<�1��<�2 ��<�	0��T��l��5J�l��cC���9�%�MCR��P�2��`�Q2@967��Q��8��9Z�2�TPB���P�2P7UA5@�o���
�5�`U���3 w���?AH�E�1��c�qAwl���A�1��512 f��1�u5Р���a5p$��56�+a��bQ5h��Ұ�1 @���pp�b[�538� xaB��|p�4�2��11/q5�p�4U5�P16 (߲�Pz��0��8�P����$�p�e5`�e5(�/�P`bbf>�X��$Z��U�5d�\� ~X�7 	  �ÿ8 k_kv��7s9 s�82 &�H5��E6���p����Ah���ñ���3J"ܫ`��4 3Ȥ59Jѧ6�0t���8��q6D0$�$�4 7���!���<�j670\tchk<�Ps0��<�B<�90��7�H<���<�\K�<�q�� ��A�C<���q�<����<�t��sg<�lc$���FA<�H��<�`��<Я���<�hk�� <Щ�B<е�o�<����<��K�<�dflr0��<Ш��� ��oҠ`���D�;�<�gEvam����B<г�o������<а�KЀ�creexl����P��<���|���j6<�s��prs.`���\���<�7������f�sgn��P�b�t�at��<�L��1B >!�svsch/  �Servo S���ule>�SVS��44�1u�_<���� (����ched���,��~��A\�� �� B���B�qA�����cj�� � 5��1<���Ә�p�css "ACS<� &(��6� �����c el���Q���~��torchms�n<�- T�Ma`�x����09 J5;�598 J681
s�7� 8��b���<Чa����te,�s�����/�E��s m��ARC.�� 1q�4�!=��C�tc�pA�@t�L��f� F����7#�2x�SE�r����UtmS�0960'���RC���`���� p��96G0= '��"H5W�� ��L���\f��� �PATb���`!40U�#!Stmt��E ��� �pMA��!p��z�2?�inA_<�X��r�X e/	cW����V���чetdl�vߏ\oveto���܏��mmonitr�0\��|#�0st��?.6a��PP����! Q�!y`�`am9e �Arol�c�43�0 �p��6��01� 25��  �<� ?v	�v	�A@�818\n; <s��I�B�2�pMPTP�"��C�1mocol��,��CT�v�'!� 0�A���8P53��y`_Touchs�s�`��<��J5���� �`mP����n[PQ �a,�E�a��IP&
&�Pth�A<�KF#R��m;�Qetth�TGHSR'�q-�Rt��o "PGIO�#�!$s�ISwka�"W�K��!�MHqH+54��5w5n/�Sm/��@ 7�*�da���8`!w/Ac��tsnf Tk�/�#gb��a��u`��^m�`u ��Zӭ�ܱQp�є� #���Ka<��M��t5QtZ�a<��dFS�5GK����G�1or��dW��64��tPx� ��P ����x,�� ?$���P<�Z4e7�g "SVGN.o�x�copy "C�O;�Wj$�O�A�9� "FSG�ѧ�%7���_��f� wQSW�F*!"(�sgatu`ɀ���_
��tp_�TPDo��9�7�9�#dߎ?���h�G�AT���!#��  �Гf�` ��" /� �w�Z� �b?6?�  ����� ���E ���M� �chrT� �K6K� �sms� �o6��~��gtdmen?3� �?��� ���mkpdtd2 ���, ���pdQ�X� ����� ����mvbkup.� �[�C�С��mku�no��prp���m�kl �4��s �n�iU��� �ldvrw���glg�4�� �p�棑��aut7�.pб�旐 �ַ������su3� �Ǜ�  �Ƿ� ���\ �6�b2X� ��&�� ���<��A4�  ��B�   946"� ��fB� �t\pa�ic\p4k94�7 ���F#���� �i�ctas���pa`���cc:�<��o������gen�� � $��F�lnp � �����stf@��1��wb�O�c��Ջ�`��߄�vri�ߢ�а�-T�� ���p�flowl� OPAc��ow���R50qtS �#T� (A��4�#���pѣV�cu3�QF�� ��SI�ac����4�6����s&��pa���!!���� ���55 �b �o)�p���0娿>
�afcal3�P߁ ��f��}���`�f��m	߳�p�d�m�/���a/��$C`ѷ��� �! track�\P� 0�ine/R?ail Tr�]T�J�69W�T  (L ��8(`љT.�`�%���D��P0� (��8�48��_ɛ�⇒A4����� �3�b13���alV@ ��NTf���%��Ii�n]0m���aen ������&?5�c@Itst3@��$� ���`�,R9�%����0氱%��pop_eners-OW �dDev��F�M�6 W���|A�Pc"�l!esv� �,��R��V$��Q���U<�V$ �k9j �6��# ������%paop/!OP�NU�V ��2celL��8g_��/�6��tscG��$���V!�3� 5vro!p�ߡ�7`�n(`� V"2D�a V'O$:S|9��� PumpE� �jQ�@�" ��!
��@бMSC#�@��)P��A�C�`��� � �v���� \mhplug�@g�"7Pb��uK")㠱io7��CJ0��E�LIOj q1g 7A93շ��5 q9 t����4.rb ST��R��CP�J989�P�LSQE�' �e C3Q(P �/Ov���o�P�� ? I1�R���5�5��f�I1`�tcm;io��MIO������Utco1"CL0�1V �cBK`io"��uM?���Sl�I0�ߢ�Eg �o���f �1tI4\onfdtI����e%�p27�Int�e�TB CoMo�o1E�R�(do5�54 (;r>Ex,p��nR##ipc�/L>��qp5���
oQ é�1�p����7/o��j�ra�pd�CDV�_��rP�֮��qp2c�nd��s �p��a �o�r`҄�S��"�c�1a�c���2kIԿ?A�pcrt���or0�qd#��"���3p+�཈D��Џ��vr2k�0���AG�.+�η�cho�;�uCp��(� �uV630� fwe P�mී�@���,`��TX�� ��d�chp "_��(	�3�����8����\p3�v����ш�9�3�1 ������low�[ͧ���chk���㳦s��s?Ө0�i�1h���2��i�w����s?1*�-0	�:�O��vr����৓0�'���PFRA�PWat?1rne@E�P�sp�& ac5� \_A�rbo#�,�a ��g��������Q=s<�ICSP+ �9_����� �q�F�A9PH51IQK93 7��HX6hQ�]PVR`S5��fPR6� iQWPR� (P^!am S�u�"��A�I0�tpprg��0���`h�@2atk932�!��E�^�^�asc "8�C��S>i�atp�"�d��@1I�
g�dsb�lfltJA�Qsable Fau�P{C!��EV0ex/!?DSB (DC��t�$�p��X 7�  �� 5��Q�t3*�~l���td9� "!0%�(5��sb9኏���\	�6#���@5��p$D@550-Ad�just PointO"tVJ�Rs�z�@䐄��!�X_�Yj�^�0\sg��4�߼}7y�\ada�"�ADJ���j�Qe�tsha<�SHAqP�sŭ'jpo�r 4�t�!��$ ��C�|�	Tk!bRPK�AR/Qiagno�stì!O!vV6�6 J`ew0�(��L���/�&krlde� ��PP���h�U b���r3�Pp<?q��DBG2C��� �X�o�1U��� ��WT`�@ip�JCM�aipper� Opv`1Se}78 (MH GF�  ;":�&##�� a�xX�֕$��388C�P����#��9.�9C�H�g##PPk�Q��8�! �_"$�"��=0%�P��A  $��_�#%0AQ�C~2� Mat.Han�dlE��!= &�pq MPLGET�0�1(�3�Tt&P�Sٰ'�B �1��B0����&p��H ��PP �'p��@�C7�PP	�TG�tD5�}m��q�Afhnd "�F_R  ���|��PP	   xT�?Q���P(Pa��TAo�����?�pmp�aO��JP ak92�5��2`@O�JRp�sQ`B2�unLHP�Tgse�GSo1�O�W�QT��v !�R�P�tp~���JRdmoan.�@��V�!ns�hYvr�QJ�g�Q�o��jY�HS~7sl�f .��pen�PDnR(R8&���ɐ823'�� ٔq���g� ���� 1��� S�� ? �c\sltQ�!|QE�P��a�r�tPg��P�� �v��"SEDG8�s0�qtdgY T��� �vP`ho�s`<`����qc�`g
�e` op�w�a@o"�ile6�H�e�ȅnR�� x�e! j517�>Ճ��J%��e�`��Q4��Q&�L�!F�J�=�o�5�z/l17���_�œ���`C0C�  ���LANG j��A���8�����gad��X�#�jp�.�0�4�Ē�ib���s�Ƒpa����&���j539.f��,Ru� Env
������3H�z�J9�����@h�Ф
Ҕ���2�a2���� (KL�n-TimФ�⠤���p�3�TS����\�kl�UTIL"�o���x�r "QM�Gl��!������1� "��S�T3�\kcmno��SФT2����ut�.�lrgeadc�}�exY�(ܤ�r��\��l��Ф�w�3��2C�*� - �C�D�E!Ĥ� .��C� R CV̴�Ҁ�C\p�Р���pďtbox��.�@�c�ycsL�:�RBT�E�veriOPTNE���;ӕ�k��e�ߦ�a�ߦ�hg��ߥ�DPN��gp�.v��r�ptl�it��0�4��te\cy����tmnu3`�r�����5UPDT��������駣��i�te �� swt�o�,���oolB �F"�Y���Q��(q��gr3��䪒��"�䴁w������߳��s��������������lS���bx " O�� ����l����0P���A�l\t�� ���������	�Colr�e!��R C��r��&r �m;`��Chang�Lq�T1 �rcm3�"��
�� 6���"����sP70���"��22!2��2D4�57�� CCF�M�H��accd	a��Q�c' ��K�@�0���K!����mo! ���,$Á��!"
 ����/�/����	Y�`,$��)�,$sk����m rC%tS1,$+�x��k1�%unc.,$poñ�1��sub��p����1��cce�5 /!&��-/?-W/i&vs�}/�%#�#�/�.@C��/� C%
�@? U ��&+��F:qt�
pD�Ѓ D	 � U�:7�Dxmov.�P��DPvc5Q.�tfr@PeC_UY?geobdtg_y[�tu���P���PTUt$�P�Sx�_�^z�_�\gvar�_�\xy�_.�[pcl`c�P���P�Ue�Pgripssuaoskuti��|�ovfinfpo}��o�j�b�P���Qud�\�aX��Pc�\Rrp��Qnƅ�P�v�P)tm�#qƆ�P�v�a+rog��a��\Q�?a+rpal?a{�{spa���P �u�Q�t�_TZp�0�osipkag3r�ovlclay(�:�t�pT�d�pu?a�c�A������KtKa�P��r��qTf|rdm���{rin#r���s � �2���|s�Pd�&v�tv��v�h�0���ystn* џ�yt'�1�p��D�p�uϑ�#�ul�@o�W6�2�siupdl�]�o�#vr�on��`1L�zp�`\�r���il3F$|l4��ǉ#q54�FyB�Տg{�`���{w�cmס���wxfe�r�UYtlk2pyp߿UYconv���sicnv�Qʯxaqg��H�Z�lct`a�o�=�p��׭nit�0믁�3������ � �� v�	�v	$��a�lϑpm�r&�B�e Wa���f�%���� ��I��߬�u�ͬ�Ka�mT�f���c��w��roǁ#�5�����?� sm��y�a��y넑 ������`����͐ϑ��p��m�Wa�1� ��A�6�S�e�X��� ��\Q}����������� ĥw߉�西߭���� ��#q0��rs�ew�@��1�a��z긱n@��.�۲;�d�������  � A�d	T$�1 pc! P��e �e� 	lf@C�@��s/�  ?�����8�� �������re�g.�C=��o�99 ~@�����$FEAT_INDEX  z ��e�� ILECOM�P :���1!!z$#�SETUP2 �;1%;"� � N f!$#_AP2BCK 1<1)?  �)��/��/  %�/�/e 4 �/�/>%�/$?�/H? �/U?~??�?1?�?�? g?�?�? O2O�?VO�? zO�OO�O?O�OcO�O 
_�O._�OR_d_�O�_ _�_�_M_�_q_oo �_<o�_`o�_mo�o%o �oIo�o�oo�o8 J�on�o��3� W�{�"��F�� j�|����/�ď֏e� �����0���T��x� �����=�ҟa���� ��,���P�b�񟆯� ����K��o����� :�ɯ^�����#��� G�ܿ�}�ϡ�6�H� ׿l�����ϝ���@)�t Px/ 2� �*.VR��߅�*�@߂�F�j�T���PCrߛ߅�FR6:����V���z�T �!���K� x��q�S�*.F�D���	�Ӑ���^�<���STM ���'���S���i�Pendant �PanelS���H I���9���U�������GIF0;���8�����JPG���;��]oR�
A�RGNAME.D)Ty�>�\"���Rc	PA�NEL1Y�%@>��e�w��2��A/�//���/�3 _/�/��/p/�/?�4�/I?�7?�/?�?�TPEINS.gXML�?>:\�?�t?�1Custom� Toolbar��?Q�PASSW�ORDg?w�FR�S:\:O�? %�Password Config{O R��OSO�O�O��_�O B_T_�Ox__�_�_=_ �_a_�_�_�_,o�_Po �_Io�oo�o9o�o�o oo�o(:�o^�o �#�G�k� ��6��Z�l���� ���ƏU��y���� ��D�ӏh���a���-� Q���������@� R��v����)�;�Я _������*���N�ݯ r������7�̿޿m� ϑ�&ϵ�ǿ\�뿀� �y϶�E���i���� ��4���X�j��ώ�� ��A�S���w���� B���f��ߊ��+��� O���������>��� ��t����'�����]� ����(��L��p ��5�Yk  �$�Z�~ ��C�g�/� 2/�V/���//�/ ?/�/�/u/
?�/.?@? �/d?�/�?�?)?�?M? �?q?�?O�?<O�?5O rOO�O%O�O�O[O�O O_&_�OJ_�On_�O _�_3_�_W_�_�_�_ "o�_FoXo�_|oo�o��o�`�$FILE�_DGBCK 1�<���`��� ( ��)
SUMMAR�Y.DG�oblM�D:�o*n`D�iag Summ�ary+8j
CONSLOG q�n�=qConsole log��7kpMEMCH�ECK��2���qMemory �Data3�;g� �{)�HADO�W(�����C�S�hadow Ch�anges���c-���)	FTP������=��qm�ment TBD�;�;g0<�)ETHERNET0��`n�q~���=qEthernet �p�figurati�on��B`%�DCSVRF/��'�@�C��%� verify allC�ޑc1p� �DI�FF8��0�ůD�{%Z�diffǯ{��q�1������J�� X�q�|�	�CHGD�&�8��ͿD�ܯ�����2pĿ����R� `�yτ�GD�.�@����D�����FY3p�ϳ���Z� h��ߌ�GD$�6�H����D�����UP?DATES.$�
�~ckFRS:\"��c�>qUpdates Listc��`{PSRBWLD'.CM��blN���e��pPS_ROBOWEL\�6o+�=� loa��o����&���J� ��n�����9��J o���"��X� |#�G�k� d�0�T��� /�C/U/�y//�/ �/>/�/b/�/�/�/-? �/Q?�/b?�??�?:? �?�?p?O�?)O;O�? _O�?�OO|O�OHO�O lO�O_�O7_�O[_m_ �O�_ _�_�_V_�_z_ o�_oEo�_io�_zo �o.o�oRo�o�o�o �oAS�ow�* ��`���+�� O��s������8�͏ ߏn����'��� �]� 쏁������F�۟j� �����5�ğY�k��� �����B����x������C�үg�v��$�FILE_N�PR�]���Y�������MDONLY 1<��~U� 
 �� ۿ(���L��5���Y� �}Ϗ�ϳ�B����� x�ߜ�1�C���g��� ��ߘ���P���t�	� ��?���c�u��� (����^������� $�M���q� �����6� ��Z�����%��I [���2��~��VISBCK��|��ų*.VD�|*� FR:\�V� Visi�on VD fileVd���� ���	/./�R/� v/�//�/;/�/_/q/ ?�/*?<?�/`?�/�? ?�?�?I?�?m?OO �?8O�?\O�?�?�O!O �O�O�O�O{O_�O!_ F_�Oj_�O�_�_/_�_�S_�_w_�_o~�MR_GRP 1=���LeC4  ;B�`	 ��lo�~li`۬B���D��fn�ӺMT� �?�� ����e`i `a�o�khb�h�o�d�cic.N���uL#2L
��|N���H�BVE��|�i`�?{��Aǿ�@i=F
��A S�8�[o�l}AĽA�߻A���s|�z�p�l}F@ �q�hq�y�~g�fF6��D�MqD��� BT��@���Ô~pD��6����l���5�?�5��|��~��� B��B��%A��B�>zBZw�~�A�B*~B�6��A��9B O7B�Bl叐�A������A�܏e�P���t����@�bo=�?��@�	Ƙ��� �Ο��+��O�:��_���p�����eBH` �Ă��a?T#=���'��d
��Z��WZ��q��Q�HZ��@����@�33@�N���\��[���ѿ��@��񿋯�*π�N�9�r�]ϖρ�<��G�=�<��m]<�+=~�m<c^���8eN7���7ѷ7�x;7;��51���	�P���?߾d2^`Yb`U�b`�����Fߪ`Үb` b`�0�����C�^o�߂o �o�߸o��o�� ]� (߁�l�������� ����#��G�2�k�V� {������������� ��1 ��-� )������� 0T?xc�� �����/')� '/M/_/q/8��/�// �/�/�/�/?#?
?G? 2?k?V?�?z?�?�?�? �?�?O�?1OOUO@O RO�OvO�O�O�O�O�� _��J����`_*�_ N�_�O�_�_�_�_o o'oMo8oqo\o�o�o �o�o�o�o�o�o7 "[Fjh�x �t��!��E�0� B�{�f�����Ï��� ҏ����A�,�e�,/ ���������/�J�� ��=�$�a�H�Z��� ������߯ʯ��� 9�$�]�H���l����� ɿ��ƿ���#��O�O V� _z�D_V_��z_�� �_���
�C�.�g� Rߋ�vߛ��߬����� 	���-��Q�<�N�� r��������� )��M�8�q�\����� ������������7 "[Fk�|�|� ���֟3�W Bg�t���� �/�///S/>/w/ b/�/�/�/�/�/�/�/ ??=?(?:?s?:�L� �?p��?�Ϧ� O��$O ��T?]OHOZO�O~O�O �O�O�O�O�O_5_ _ Y_D_}_h_�_�_�_�_ �_�_�_o��@o
�go *owo�o�o�o�o�o�o 	�o-*cN� r������� )�;�M������� ��ˏݏď��%�� I�4�F��j�����ǟ ���֟��!��E�0� i�T���x���ï�?�? ��O��?OO�t� >O������ѿ��ο� �+��O�:�s�^σ� �ϔ��ϸ������ � 9�$�6�o�6o��Zo�� R����������5� � Y�D�}�h������ �������
�C�U�� y�����d�����:��� ��+Q8u` ������� ;&_Jo�� ����//گ4/ ��x�j/4��/X�n/|� �/��/�/!??E?0? B?{?f?�?�?�?�?�? �?�?OOAO,OeOPO �OtO�O�O���O�O_ �O+__O_:___�_p_ �_�_�_�_�_�_o o oKo6oooZo�oZ��o �o�o�o��xo
G 2kR����� ����1��.�g� R���v�����ӏ��� 	��-��Q�/*/�� N/��r/�/ޟ�/��/ )�D�M�8�q�\����� �������گ���7� "�[�F�k���|����� ٿĿ���O�O�O��W� B�{�fϟϊ��Ϯ��� ������A�,�e�P� ��t߆߿ߪ��ߪo� �+�=�a��߅�p� ����������� � 9�$�]�H���l����� ����������#G�2W}h�p��$�FNO �������
F0� �  >#�1 D|�� �RM_CHKTY/P  � �q�� ��� ��OM�� _MIN� m�����  X�� SSB_CFG� >� ~�Jl�Aj�|�TP_DEF�_OW  m�|��IRCOM� ���$GENOV�RD_DO�ܠ��THR dz�d�_ENB�� �RAVC_?GRP 1?3� X�e/��/�/ �/�/�/�/�/�/? ? =?$?6?s?Z?�?~?�? �?�?�?�?O'OOKO 2OoO�OhO�O�O�O�O��O�O�ROU? E\� q���|���8�?#��O__K_m_o_ꐖ  D3���_E�_2q�@A��\Bȡ��Rp��>Y_6 SMT<#FC-�Ufoxo�o��HOSTC,1G�Y?��_ 	��h�k�o�f�oyeCUg y�z1�������p	anonymous�5�G�Y� k�w��o�o�o��� ���*�<��`�r� ������ˏ	���� �&�8����������� ���ȯگ���M�� 4�F�X�j�����ݟ�� Ŀֿ���I�[�m�� ��fϵ��ϜϮ����� }�����,�O�Pߟ� t߆ߘߪ߼���/� A�C�(�w�L�^�p�� ���ϸ���������� a�6�H�Z�l�~����� ������9� 2 DV��z���� ��#��
.@�� ������������ �//g</N/`/r/ �/����/�/�/? Qcu��/[?��? �?�?�?�?)/�?O"O 4OFOi?�/�/�O�O�O��O9m�aENT 1=H[ P!^O_  `_?_._ c_&_�_J_�_n_�_�_ �_o�_)o�_Mooqo 4o�oXojo�o�o�o�o �o7�om0� T�x����� 3��W��{�>���b� ��Տ���������A� �e�(�:���^������㟦�QUICCA0�̟ޟ?��1@��.����2��l�~��߯!ROUTE�R௼�ί/�!P�CJOG0��!�192.168�.0.10	��GN�AME !�J!?ROBOT���N�S_CFG 1G��I ��Auto-sta�rted/4FTP:?�Q?SOBχ? f�xϊϜϮ��?���� ���+�߿�P�b�t� �ߘ�6�����(� J� �1�C�U�g�6ߋ� ���������x�	�� -�?�Q�c� ?2?D?�� �������)�� M_q����:� ��%t����� m�������� ��!/3/E/W/z{/ /�/�/�/�/�/6H Z ?n/S?�w?�?�? �?�?�/�?�?OO<? =O�?aOsO�O�O�O�/ 
??.?0O_d?9_K_ ]_o_�_PO�_�_�_�_ �O�_�_#o5oGoYoko �O�O�O�O�_�o&_�o 1Cogy� ���oT��	�� -�|o�o�o�o����o ��Ϗ����)�;� M�_�q��������˟�ݟ�ÿT_ERR� I�����PDUSIZ  ^���$�>=�W�RD ?޵w���  guest+�}��������ůׯ��SCD_GROUP 2J�W �`�1���!��L_��� � ��!�	 i-y	�E���Q��E EATSWI�LIBk�+��ST� 4�@좰1��L�FRS�:аTTP_AU�TH 1K�<!�iPendan�������!KAREL:*���	�KC�.�@���VISION SET���u���!�ϣ��������	� �P�'�9߆�]�o޽�CTRL L���؃�
��?FFF9E3��u����DEFAUL�T��FANU�C Web Se/rver��
��e� w���j�|��������WR_CONF�IG MY��X����IDL_CPU_PC����B�x�6��BH�MIN'��;�?GNR_IO�K����"��NPT_S_IM_DOl�v��TPMODNTO�Ll� ��_PRT�Y��6��OLNK 1N�ذ��� 2DVh��MA�STEk�s�w�O>ñO_CFG��	�UO����CYC�LE���_AS�G 1O��ձ
 j+=Oas� ������//\r�NUMJ� �<J�� IPCH�x���RTRY_CN��n� ��SCRNO_UPDJ����$�1 �� �P�A���/���$J23_DSP_EN~���p�� OBPR�OC�#���	JOGv�1Q� @��d8�?� +�S? /?)3POSR�E?y�KANJI�_� Kl��3��#R������5�?�5CL�_LF�;"^/�0EY�LOGGIN� �q��K1$��$L�ANGUAGE YX�6�� vA��LG�"S�߀������x��i��@Z<𬄐'0u8������MC:\RSCH\00\���S@N_DISP T�t�w�K�I��gLOC��-�DzU��AzCOGBOOK U	L0��d���d�d��PXY�_�_ �_�_�_ nmh%i��	kU�Yr�Uho�zohS_BUFF [1V��|o2s� �o�R���oq��o�o# ,YPb��� �������(��U��D/0DCS }Xu] =���"l ao����ˏݏ�3n��IO 1Y	 �/,����,�<�N� `�t���������̟ޟ ���&�8�L�\�n����������ȯܯ�E�e�TM  [d �(�:�L�^�p����� ����ʿܿ� ��$� 6�H�Z�l�~ϐϢύdN�SEV� ]�TYP�$���)߄m�1RSK�!O�c>�"FL 1Z�� ����߯������ߘ��	�:�TP5@����A]NGNAMp�$�E��k�UPS P�GI|%�1�%x�_�LOAD0G =%Z%TEQѼ���MAXUALRM;'�I(��~���#�� V�#a��CQ[�x�8��n��"�1060\.	 �F�	�Ϣ� ������������  D'9ze��� �����R =va����� ���*//N/9/r/ �/g/�/�/�/�/�/? �/&??J?\???�?k? �?�?�?�?�?�?�?"O 4OOXOCO|O_OqO�O �O�O�O�O_�O0__ T_7_I_�_u_�_�_�_��_�_o�_,o��D_LDXDISAc����MEMO_A�P]�E ?��
 �5i�o�o�o��o�o�o�o��IS�C 1]�� � oTd��\no� �������� I�4�m��f���$��� ������!��E�Ə T�f�:�����ß��� ��z��ܟA�,�e�w� ^������~����� � �=���L�^�2��� ������߿�r� �Կ�9�$�]�o�(t_MS�TR ^�͂�S_CD 1_xm�W� ��S�������=�(� :�s�^ߗ߂߻ߦ��� ����� �9�$�]�H� ��l���������� ��#��G�2�W�}�h� �������������� 
C.gR�v� ����	�- Q<u`r��� ���//'/M/8/ q/\/�/�/�/�/�/s��MKCFG `���/��LTAR�M_2a��2 �#\`Y>G`�METPUT`�"�����NDSP_CMNTs506�5N�� b���>�"�1�?�4�5POSC�F�7�>PRPM��?�8PSTOL �1c2}4@p<#�
aA�!aEqOG]O O�O�O�O�O�O_�O �OA_#_5_w_Y_k_�_��_�_�_�Q�1SIN�G_CHK  ~+O$MODAQ73�d
?�7:eDEV� 	��	MC}:MlHSIZEs0����eTASK �%��%$123456789 �o��egTRIG 1�e�� l��%��?   A$��F�fYP�a,u��c�EM_INF 1�f>7 �`)AT&FVg0E0N�})�q�E0V1&A3&�B1&D2&S0�&C1S0=�})�ATZ�� �H@�E��q9m��xAu�@��X�������� � �����v�)��� я��П�������*� �N�����7�I�[� ̯ן���9�&��� \����g�����i�ڿ ������ï4��XϏ� iώ�A���m������� ߿�ѿB����ϊ� ��O������ߟߩ�� ��>�%�b�t�'ߘ�K� ]�o߁�����(�_� L���p�+���������~�.ONITOR�0�G ?ak   	EXEC1�#�2345��`789�#��xx x*x6xBxN�xZxfxrx2�2�2�2�2��2�2�2�2��2�33�3�aR_GRP_�SV 1g�y�a(��Q>`�?��뿲��cj��?�ZF@K�	Hm�a_Di�n�!�PL_NAME �!�5
 �!�Default �Personal�ity (fro�m FD) �$R�R2� 1h)d?eX)dh�
!�1X d�/d/v/�/�/ �/�/�/�/�/??*? <?N?`?r?�?�?�?�?�?�82S/�?O O2O�DOVOhOzO�O�Ob< �?�O�O�O�O_"_4_@F_X_j_|_�_LhR�g 1m)9`\bO0 �_pb�Q� @D�  �Q?���S�Q?`�QaAI�Ez  a�@og;�	l�R	� 0`4b@(4c.a�P�Jd�Jd��Ki�K��J���J���J�4�J~��`jEa�o-a�@��o��l[`@�z�b�?f�@�S��a�Q��o�c�=�N���
�����T/;f��`��l[`��*  �p  ��$p> p�$p���o?p?����{�����o�Bntr�Q�skse�}�l�p�  ��pu`j  #p��vks��� 	'� �� �I� ��  ���}:��È6�È=��9�N��b@^�d� �n�Q���{�R�x���nN. ��  '����a�`@a�@��t�@p@p@�CpC0�fT0�+pB/pC3}�PO�@%�Eab�oo$|m�����gA %���. ���z�`�P���QDe���˟���(��m�� ��t O� �ru �4 ��R�c��s� :��u�a�P�` �?�ffb�!�����>7� ��گ�0�af��>搠���iP�P;�e�S�Ea4f�u�>LX��s�b�<	�I<g��<#�
<2���<D��<��
0vo��¯�S��S.����?fff?u�?y&찗d@T����?�`?Uȩ?X����Z�� �T:z�TB��Wa�з*d ů�ρϺϥ�����߀��&�8�#�\�h�+�F. Kߘ�G߼�3����Wɯ���G�@ G����X�C�|� g�y���������j Z���ￏQ����� ������3����� ��/A��t_������������b���@+FpؠIP�t��%���[`B�0�����<ze�cb!@I��
�M`B@���@`�9@y���?�h� ��@�3�[N���N�N�E���<�/:/L ��>��ڟ�A��p�C�F@��S�b/DpX������@�t���%�h��`/qG���GknF�&�FצpE�,8{�/ F���ZG���F��nE�DE,�ڏ�/� ���G���F7��F?��ED��.�� C?.?g?R?d?�?�?�? �?�?�?	O�?O?O*O cONO�OrO�O�O�O�O �O_�O)__M_8_q_ \_�_�_�_�_�_�_�_ o�_7o"o4omoXo�o |o�o�o�o�o�o�o 3WB{f�� �������A� ,�Q�w�b��������� �Ώ���=�(�a��L���p�����(r!3g�ji��r������3Ա�ڟ�y��4 ����y���P�2�D�&�j�b^�p�1w���������ʯ���Pܯ� �s�P^�PD�c�`�m���y�\������Ӱ�¿Կ��� ��.�G����}� �ϡ���홍�U�_�J���$�y.�@�v�d� z߈ߚ�x�4�����ߠ�� ��D�.�2� ��$[�G�[�^�Bh���B��CH�  ^����u�����������p�h�M�_�q�P���������^��^�Y�m�2��
 ����#5G Yk}�������h*�� ��>�x�}��$MSK�CFMAP  ���� �����m�N"ONR�EL  6��9_�"EXCFE�NBk
7]�F�NC�}JOGO/VLIMkduy]d"KEYk�]"RUN���"SFSPDT�YU��v_SIG�Nk}T1MOT��z"_CE_�GRP 1n��9\���/���/�/ 4��/?�/2?�/'?h? ?�?C?�?�?y?�?�? �?O�?@ORO	OvO-O oO�OcO�O�O�O_�O�*_<_#_`_-�"TC�OM_CFG 1�o/���_�_�_
�|Q_ARC_��6��UAP_CP�L�_�NOCHE�CK ?/ 5�;h9oKo]ooo �o�o�o�o�o�o�o�o�#5GTNO_?WAIT_LF'56y"NT�Qp/����q_ERR�!29q/_�� R_���"�:�L�d�T_MO�sr�},� #<P_��_�P�ARAM�rs/������MW���� =e�345678901.�@�R�)� q���_�����˟����ݛLW�3�E�؏�i�cUM_RSP�ACE,�������$ODRDSP�S�I&�OFFSET�_CARToݨD�IS�ݢPEN_FILE�I!�Q�v��POPTION_�IO���PWOR�K t�'� QT�|�
� ^�F�� �
���Z���	 �m���A�
��i��_DSBL  Ķ�v���ޡRI_ENTTOj��C���8�ῠUT�_SIM_DJ��6	��VàLCT u�}\��Q��>W�_PEXE���RAT���� ��>�UP ve�����������*�8���$��2�#h)d�eX)dh�O�X dY�ߑߣ� �����������!�3� E�W�i�{������������2n��)�;� M�_�q���������<�����+= Oas���X���� O��1m(��O�(�.�g��"0 �дu� � @D�  �?���?рH�D4  EzZ3�;�	l	 '0ӀS@SM�� �i�i �H)�!H,�H�8�Hm�G�?	{G�8��6��MV��� �C�)���)�����Ճ�*  �p W � > � p,�//)/ B,��Btr�«��H�¼�/�� �/�"�# �,0 ��� �  z� ߽pj  B ���&X�?MU	'�� � 12I�� �  �=��-=���U?g;/�@}?�0~.ѱ��?;Ѳ���H[N5��?  'M�D��> C)�f)�J B�N +��=%O7O�R��@D1�oo�$����JWAD0�J5�4�: �1�E&?��O�O#__G_2]��� �t O�� ru �4 ��R�UɳO� :�%Ёр~� �?�ff��@[�_�_V_{�o~�b�18р"o0j>�P�Q6YPрZo�WrAd<S�%�>Lw0�#��<	�I<g��<#�
<2���<D��<��`��l�_�ѳ|Mb�@?fff?�0�?&p:T@T��q?�`?U��?X�-q�iyB q5Ya��g I�_������ !��E�W�B�{���d� ����ՏLnpΏ/�~ʈG�@ G�� U�ȏy�d�������ӟ �������yB=� � �?p���/򏸯�߯ R���'�9��oN�`������~�����ۿƿ�B�ĮD�e�ֿ;�xҿ_�J�?��h�PoϨϓϸ��D4��b!�_@���� ߧ�������%�@I��)�M`B@���@`�9@y���?�h	� ��@�3�[N���N�N�E��<��/Y�kЖ>���ڟ�A�p��C�F@�S����pX������@�t��%��h��߉!G���GknF&��FצpE,8�{�� F�Z�G���F�n�E�DE,ڏ���ૐ�G���F7��F��ED��Mf��b�M� ��q��������� ��(��8�^�I���m� ��������������$ H3lW�{� �����2 VAS�w��� ���/.//R/=/ v/a/�/�/�/�/�/�/ �/??<?'?`?K?p? �?�?�?�?�?�?O�? &OO#O\OGO�OkO�O�O�O�N(]�3�j�i�O�a��	U�E3�Ա��O_<q4 ��%_7_<q�Pq�Q_c_ERjb}_��_1w������]�Y�_�_o�_1o�l��P�bPcn~� ��o�O�o{_�o�oY�`��o�o,/; M#�f0o���� �Y�et�~�i#�1�C�yM�_��������� ��{bS�Ԏ��	�?�h-�c�Mj2���$�V'G�z}�B����B��CH�}�9� ֟�����0�B���wl�~�������Ư*�T���\�r�qQ��U
 ί �0�B�T�f�x����� ����ҿ���χ���� ��]{x}���$PARAM_MENU ?Յ��  �DEFPU�LSE�	WAITTMOUTl��RCV� �SHELL_WR�K.$CUR_S�TYLj���OsPT����PTB�����C��R_DECSNw�Te'�!�3�E� n�i�{ߍ߶߱������������F�A�US�E_PROG �%P�%B��V�CC�R��UeXÚ�_H�OST !P�!�����Tt`����Ŀ�����4���_T�IME�� �T�  �A�GDEBUG���P�V�GINP_�FLMSK]���T�R����PGA�� 2|�[���CH�����TYPEM�Y� A�;�Qzu��� ���
)R M_q����� ��/*/%/7/I/r/ m//�/�/�/�/�/?���WORD ?	>��	RS��C/PNS�E��>2sJO���BTE����TRACECT�L�PՅZ� }{`� a`�{`�>q6DT QexՅ�0�0D���Sc{aa�0���2���?T�?�2�4D�2#A�O.O@ORF�cA�bB`D	`D
�`D`D`D`D�`D`D`D`DB`DObOtO�F A �5P�2Q0TOBPR PBP�BP0T�B@P�BP�BP�A,_ >Z�_=_O_a_s^$_�_ �_
b��"o4d�_�_�_��O�O__a�1	a�d�TVd^dbfdnb�Wr�k@}�o�o�j;qwc�TvT~T5OcM_ q�����v,> �
�t�@�R�d�v� ��������+���� ��ˏ��,�>�P�̟ ޟ���9�*�<�N� `�r���������̯ޯ ���&�8�J�\�n� ��������ȿڿ��� �"�4�F�X�j�|ώ� �ϲ����������� 0�B�T�f�xߊߜ߮� ����������,�>� P�b�t������� ������(�:�L�^� p���������������  $6�Fl~ �������  2DVhz�� �����
//./ @/R/d/v/�/�/�/�/ �/�/�/??*?<?N? `?r?�?�?�?�?�?�? �?OO&O8OJO\OnO �O�O�O�O�O�O�O�O _"_4_F_X_j_|_�_ �_�_�_�_�_�_oo 0oBoTofoxoN�o�o �o�o�o�o,> Pbt����� ����(�:�L�^� p���������ʏ܏�  ��$�6�H�Z�l�~� ������Ɵ؟����  �2�D�V�h�z����� ��¯ԯ���
��.� @�R�d�v��������� п�����*�<�Nπ`�rτϖϨϺ�����$PGTRACE�LEN  �� � ��������_UP _y�����������_CFoG z��������<��� �<�Z�l�<�$�DEF�SPD {/�l�a�����IN'�?TRL |/�S��8Lԃ�IPE_C�ONFI+�}�O��<�x�WLID(�~/��?GRP 1���������@�
=��[���A?C��C
�XC)���B��r������dL�z������?� 	 r�N�8�Ҩ�� ´�����B������������A���> �6>�7�D_������� �='�=)�� ��������	B-���Q�M��� G Dz����
� �&L7p[� �����/��6/!/Z/��
V7�.10beta1�<�� B=q��"`ff@��"�>����!=�̽͏!A>ff�!@w�ff�"�\)�"D��?�  �!1@�!� �!Ap�#W��h/??*?<?K;�w����O/�?K/ �?�?�?�?O�?O>O )ObOMO�OqO�O�O�O �O�O_�O(__L_7_ p_[_m_�_�_�_��_  o�_$oo!oZoEo~o io�o�o�o�o�o�o�o� DQy{/�#F@ {yw}�y{ջy �-������/�Z? l?~?w���t�����я ���������O�:� s�^���������ߟ� ܟ� �9�$�]�H��� l�~����_ۯ��� ��5� �2�k�V���z� ����׿¿�����1� \n�j�|϶�� �����	�4�F�X�j� c�χߙ߄߽ߨ��� �����)��&�_�J� ��n��������� ��%��I�4�m�X��� ��ί����������! E0B{f�� ����H�Z� ��Vh�ϴϊ�� ��� �2�D�V�O/� s/^/�/�/�/�/�/�/ �/? ?9?$?6?o?Z? �?~?�?�?�?�?�?O �?5O OYODO}O�O�� �O�OtO�O�O_�O1_ _U_@_R_�_v_�_�_ �_�_�_"4FxBo |����o��o�o //0/B/;�__J �n������ �%��I�4�F��j� ����Ǐ���֏�!� �E�0�i��O^���N� ß՟�������A� ,�e�P�b��������� �o o2oTo.�hozo �o�����o��Ϳ�o
 گ'�֯K�6�o�Z� ��~Ϸ��ϴ������ ��5� �Y�D�Vߏ�z� �ߞ����������1� �Uy��:��� ������	���-��Q� <�u�`�r��������� ��T�f�x�n ��������� ���7"[Fj �������!/ /E/0/i/T/f/�/�/ �/�/�/�/?�//?A? l�e?w?&?�?�?�?�? �?�?�?OO=O(OaO LO�OpO�O�O����* �O_@RdZ_l_���$PLID_K�NOW_M  ~���A��TSV ��]�P�[? �_�_o�O&oo#o\o��B��SM_GRP� 1��Z� dI`~�oo$Cf~�d����D��TPbj�oLk�f�o "~�U�o>n2 T�~����� 7�4���p�D���R� ��ʏ����������6��
�T��*������QMR�c��mT�EGQK? GR��(�#��� [��/�A�S������� �����$����W�� +�=�O������������� ���S�Ͻ�S�T�a1 1��ڗ���P0� @����E�ϲ������ ���M�0�B�T�fߧ� �ߜ�����������7�P�,�m��2����N�A�<��z�3��������4���������5)�;�M�_���A6x���������7����������8(:�L��MAD  ����� ��PAR�NUM  ���Ko���SCH�
 ��
��S+UPD��xaq{��_CMP_�`� <P�z '�U�ER_wCHK����Z���RS���_�QG_MO� �%_�~�_RES_G����� ��v/{/�/ �/�/�/�/�/�/*?? N?A?r?e?w?J'��W,g/�?L%��?�?�? N#(��?OON#w�4O SOXON#��sO�O�ON#  �O�O�ON#d �O_<_N"V 1��Uua^�@cX��Pp�P_$@cW،P��P_@@cV��P�"THR_INR���pbA%d�VMASmS�_ Z�WMN�_��SMON_QUEUE ��e��`UȨ`�N�U�qN�V�2`END4a6/NiEXE]oNeW�BE\`>o/cOPT�IO;g?+2`PROGRAM %j�%1`O_�0bTA�SK_I��nOCFG �o�^9pDATAɓ�B{@ev2w��� ���z��+�=�O���s���������nzIWNFOɓ��}�!d r��!�3�E�W�i�{� ������ß՟���� �/�A�S�e�w�҇ބ���| �98q�DIT �Bׯj~WERFL~hwS~��RGADJ �^ƪA�  ,�?E��8��Q�IORIT�Y�W���MPD�SP�a�j�U�W�vT�OG��_TGp���Rj��TOE�P�1�ƫ (!�AF�PE5 ����!tcp��%��!ud�?�!�icm<�Q_��XYm_<q�Ƭ�Oq)� *������Op������������ <�#�5�r�Yߖ�}ߺ�@�߳������&�*�OPORT�a�Op�A%�_CAR�TREP~`Ʈ��S�KSTA�X!*SS�AV`�ƪ	2500H809u�PT毙䕣�ƫ�����`X#�$�6�^m�URGEU`B��6A)WFP�DO�V�2��W�q�?Q�WR�UP_DELAY� �Ưe�R_HOT�hwR%z�����R_NORMAL��n��6SEMI�:y�QSKI�P���X%�x 	������� �X%-;%[m E������ �!//E/W/i///y/ �/�/�/�/�/�/?�/ ?A?S?e?+?�?w?�? �?�?�?�?O�?+O=O�OO1U�$RBTI�F��NaRCVTM쒻���m@DCRڕ���A@��u�B��rA��U���@�-�)�����һ;�/ž؞~����_��_ <�	�I<g�<�#�
<2��<D��<��
+_ _{_�_)`���_�_�_ �_�_ oo$o6oHoZo lo~oi_�o�o�o�o�o �o�o DV�_z �������
� �.�@�R�=v�a��� ��������׏�*� mN�`�r��������� ̟ޟ�����8�J� 5�n�Y���}���ȯ�� ���A�"�4�F�X�j� |�������Ŀֿ�ӯ ���0�B�-�f�Qϊ� m����������� ,�>�P�b�t߆ߘߪ� �ߧ��������(�:� %�^�A����ϸ��� ���� ��$�6�H�Z� l�~���{�������� ���� 2Vh�� �������
 .@R=O�s �����/�*/ </`/r/�/�/�/�/ �/�/�/??&?28�A�GN_ATC 1���K AT&FV0E02;�ATDP/6�/9/2/9p8�ATA2>,�AT%G1%B9�60k9+++��?,�1H�?,�AI�O_TYPE  �EC/4?RE�FPOS1 1�> K x�O[H/O/�O�MNO`O �O�O�O_�OC_�Og_�_d_�_+K2 1� KLON_�_o�_*o<�_5A3 1��_�_��_ o�o�o�o@oS4 1�Woio{o�o3�W�oS5 1� �o�oJ���jS6 1������]�H����S7 1��(�:�t��ݏ|���S8 1������Ϗ	���r���)�SMASK 1� O�  
���ɗXN	O�?���1.�8�1A?MOTE  �.D�N�_CFG ��U���5�0BPL_R�ANGQ�K!Y�PO�WER �Q5� a�SM_DRY�PRG %�%�R���ȥTART �����UME_�PROׯ�d�.D_�EXEC_ENB�  �5]�GSP�D=����Y3��TD�B����RMÿ��MKT_ѐT��S�D0�OBOT_NAM/E �S�;9�OB_ORD_N_UM ?��A�H80�0|I$�	��s	��\����� ���e��	@�}�D�|��D0PC_TI�MEOUT�� x�D0S232n�1��Q; LTE�ACH PENDcAN��j�5��=�Q�x0Maint�enance CGonsK"-��"+�~t4KCL/C��}�6��|� No Use�=p[߹�F���NPO��\��5�_���oCH_L@��U�曑	J��MAVGAIL`���+��]��I�SPACE1 ;2�=L  ����p��扢J@��>��8�?���  ���V�w�N����� ����������4�& G
l�}d	Q5U1� ��������`4& G
l}d�#��2�������� 2A/b/%/w/�//�/�3����	/ �/-/O/^??B?�?�?�?�?�4�/�/?? &?�?J?l?{O�O_O�O�O�O�O�5�?OO 1OCO�OgO�O�_�_|_ �_�_�_o�6_*_ <_N_`_o�_�_�o�o@�o�o�o!�75o GoYoko}o+�o�o�����)��>��8 Rdv��H��� ��ӏ%�F�-�[���G �� tR�;�
�� �� ��ԟ���
��.�@� ���c���p���8�¯=�dؠ��ϟ���!� 3�E�W�i�_�q���� ��x��կ��'�9� K�]�oρ�w��ϛ��� Ͽѿ����5�G�Y� k�}ߏߡߗ��߻������� `S� @��8堯F�"�*ل�����߇�� �����,����V�h� 2�<�N����������� ��.L4v��R\n�����
�f�7�_MODE�  ��MS E���&����Ïb��*	�&/�$�CWORK_AD�]	3��!R  ���t +/^ _INTVAL]����hR_OPT�ION�& h��$SCAN_T�IM\.�h�!R� �(�30(��L8/������!��3��1��/@>.?���"S22�41�9d�4�1"3��@���?�?��?���IP���@���JO\OnOE@D���O�O�O �O�O�O__(_:_L_8O���4X_�_�_��8�1��;��o�� 1��pc]�t��Di�|1��  � lS2 ��15 17oIo[omo o�o�o�o�o�o�o�o !3EWi{� ���wc���	� �-�?�Q�c�u����� ����Ϗ����)� ;�M�_���`[���� ğ֟�����0�B� T�f�x���������ү������$�7�  0��� om������ ��ǿٿ����!�3� E�W�i�{ύϟϱ��� ����v���/�A�S� e�w߉ߛ߭߿����� ����+�=�O�a�s� �����ߖ����� � �$�6�H�Z�l�~��� ������������ `2DVP�\�  �A ������� %7I[m��������/ �/C(/N/`/r/ �/�/�/�/�/�/�/?�F;/?B?F��x1 ;?w=	�12345678�{��l�@�P�?�?�?�?�?O9/2ODOVOhOzO �O�O�O�O�O�O-/
_ _._@_R_d_v_�_�_ �_�_�_�O�_oo*o <oNo`oro�o�o�o�o �_�o�o&8J \n���o��� ���"�4�F�X�j� |������ď֏��� ��0�B�T�f����� ������ҟ����� ,�>�m�b�t������� ��ί����(��6yI�[�@�`����������Cz  B}p*   ����254F��$SCR�_GRP 1�(��e@(�l���0@} `1 [1�s	 )�3�C�<�t�vr�Y�8P�}�kϤ���[�95C����-�u��ȡ���L�R Mate 2�00iC �190��1Շ0LR2CA �3�=OÆ�D�
f؜1u�2�U7��`1��v��@�u���	t���������$�^0�2���_2T� gϡϊ��o�F�D�f?@��s�����￶ht _,Z�qO� LN�B�˰�P�N�g�N�9Aܰv�  @DЎ�rN�@����  ?� ���J�H˰��y�N�F?@ F�`���� ��A,Qwb ���n�N����0���B�� _J�n���� �/�%//I/��E+@:3��6?|?�5��
�/��/�#��@=��a"�/pǢ� 3B�07�590@7����EL_DEFAU�LT  I����� ^1M�IPOWERFL�  V�v5]2�0W3FDE�m4 v5 ��ERVENT 1O���O�t3C��L!DUM_E�IP?�8�j!?AF_INEj0O��$!FT�?=N�OaO!Q�O ��PO�O!RPC_OMAIN�O�H��O��O�CVIS�O�I���OE_!TP8PP�U<_�9d4_�_!
�PMON_PROXY�_�6e�_�_XR�_�=f�_)o!R?DM_SRV*o�99gouo!RR8�o��4hdo�o!
�@M��_�<i�o!R�LSYNC4y�8�oY!ROS�?�|�4H�tO� 8c�����;�� _�&���J���n����� �ȏڏ7�I��m��4���X����7ICE�_KL ?%�;� (%SVCPRG1�����!�"�3*�/��4R�W�"�5z���6�����7ʯϯ�C��5�	9��oG�� ��o������D��� �l��񑔯�񑼯 7���_������ 4����]�������� ���'��տO���� w��%ϟ��M���� u����������?� A��Ͽ�ђ�؟ꐊ� ��ɱ��������?� *�c�N����������� ������);_ J�n����� �%I4mX �|�����/ �3//W/i/T/�/x/ �/�/�/�/�/�/?/?�?S?Ś_DEV ��9�MC�:[8�im4O�UT_Rf1~6i8REC 1���f0�0� �1 	  �2�?�1���3OMO�@O+OdO��
 �Z����6 s + UEBf0K�q�0�0�f0ʬ��2�3%f0nf0�@ ��-�)X�O�2E0��0'qE0_�O_�5"_�C &_L_:_p_^_�_�_�_ �_�_�_�_o o"oHo 6oloNo`o�o�o�o�o �o�o D2T Vh������ ��
�@�.�P�v�X� ������Џ����� *��N�<�r�`����� ��̟��ܟޟ�&�� J�8�n���b�����ȯ ��دگ�"��3~A� (��P���t�����ο �¿��(��8�:� Lς�dϒϸϦ�����  ���$�6��Z�H�~� lߎߴߢ��ߺ���� ��2� �V�D�z��n� ���������
���.� @�"�d�R���v����� ��������<* `N��x��� ��8HJ \������G�5oV 1��< P_��1�GFO�2  �jH�0wXJa?_�TYPE�?k2HE�LL_CFG i�z:f2/ �B��/�/ %RSR �/�/�/?
?C?.?g? R?�?v?�?�?�?�?�?�	O�?-O?O/�  �!�@oO�O�O�C�I�AP�O�B�@S�WgB2Pd�O|�O�&HK 1��+ �OE_@_R_d_ �_�_�_�_�_�_�_�_ oo*o<oeo`oro�o�a&�#OMM ���/�o�"FTOV_�ENBr$!}*OW_REG_UI�o~e"IMWAIT�b��I${OUTv�$&yTIMu���`VAL5's_�UNIT�c�v})M�ON_ALIAS� ?e�i ( he!� ��$�6� Q&�c�u�����D��� Ϗ�����)�;�M� _�q��������˟ݟ ����%�7��H�m� �����N�ǯٯ��� ���3�E�W�i�{�&� ����ÿտ習��� /�A��e�wωϛϭ� X�����������=� O�a�s߅�0ߩ߻��� �ߊ����'�9�K��� o�����b����� ���#���G�Y�k�}� ��:����������� 1CU y�� ��l��	- �Qcu�2�� ����/)/;/M/ _/
/�/�/�/�/�/v/ �/??%?7?�/[?m? ?�?<?�?�?�?�?�? �?!O3OEOWOiOO�O �O�O�O�O�O�O__ /_�O@_e_w_�_�_F_ �_�_�_�_o�_+o=o Ooaosoo�o�o�o�o �o�o'9�o] o���P�������s�$SMO�N_DEFPRO ���:�� *�SYSTEM* � �l�*�RECALL ?}:�� ( �}5x�copy fr:�\*.* vir�t:\tmpba�ck��=>lap�top-u9nq�dgeh:592�8 ��3 723� 5�͏ߏ�s}6z�a��������B�T���:{�s:ord�erfil.da�t������ӟ�}=1{�mdb:��� ����=�O�a��y�� �����ү������� -�>�P�b�u������ ��ο�����)��� L�^�q�����9��� ������%���H�Z� m����5������ ����!ϳ�D�V�i�{� ߟ�1�����g��ϊ����/�@�R�d� }
�xyzrate 61 ��)�;��������!z���39020 ����?Qc���tpdisc 0,������tpconn 0 ����J\��;zߌ߂6����2�ߕ �>/P/b/�����1/�/�/g/7��/�/ �/D?V?i{�? �/�?�?g?��?/�? @OROdOw/
?O�/�O �O�O�/�O�O+?<_N_ `_s?�?O�?;_�_�_ �?_�_'O�_Jo\ooO �O_�O7o�o�o�O�O �o#_�oFXk�}��!3������7068�=�O�a��t�{b�soutpu�t\calpr.�pc�P: ove�r =>3355�4432:1000172�ÏՏh^=3z�temp���@���?�Q�c�vP4z�test.ls�� ��/���ҟ�wU����tp~��������H� Z�m��,���ϯ ���������M�_� r_�_o�6�ǿٿ�_ �_�����>�P�b�o���$SNPX_A�SG 1�������� �P'%R[1]@1.1f�l�?�o�%���Ͽ�  �����6��@�l�O� ��s߅��ߩ�������  ���V�9�`��o� ������������� @�#�5�v�Y������� ��������< `CU�y��� ���&	0\? �cu����� /�/F/)/P/|/_/ �/�/�/�/�/�/?�/ 0??%?f?I?p?�?? �?�?�?�?�? O,OO PO3OEO�OiO�O�O�O �O�O�O_�O _L_/_ p_S_e_�_�_�_�_�_  o�_�_6oo@oloOo �oso�o�o�o�o�o�o  V9`�o �������� @�#�5�v�Y������� Џ��ŏ���<�� `�C�U���y���̟�� �ӟ�&�	�0�\�?� ��c�u��������ϯ ���F�)�P�|�_��x�PARAM ���� ��	���P���p�OFT_KB_?CFG  �����״PIN_SIM  ��̶�/��A�ϰx�RVQST_P_DSB�̲�}Ϻ���SR ��	�� & TE�ST V�����ԶTOP_ON_�ERR  ������PTN z	��A���RING_PRM��� ��VDT_?GRP 1�����  	з��b�t� �ߘߪ߼�������� +�(�:�L�^�p��� ��������� ��$� 6�H�Z�l�~������� �������� 2D V}z����� ��
C@Rd v������	/ //*/</N/`/r/�/ �/�/�/�/�/�/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4O [OXOjO|O�O�O�O�O �O�O�O!__0_B_T_ f_x_�_�_�_�_�_�_ �_oo,o>oPoboto �o�o�o�o�o�o�o (:Lsp�� ����� ��9��6�׳VPRG_CoOUNT��ќ��d�ENB/�_�M���鴖�_UPD �1�	�8  
 M�������-�(�:� L�u�p���������ʟ ܟ� ��$�M�H�Z� l���������ݯد� ��%� �2�D�m�h�z� ������¿Կ����
� �E�@�R�dύψϚ� ������������*� <�e�`�r߄߭ߨߺ��������\�YSDE�BUGn�Ӏ���d���"�SP_PAS�Sn�B?4�LOoG �΅�������
�  ������
MC:\x`��a�_MPCf�΅����ҁ��� �ҁ��SAV �bi���������SV�TEM_T�IME 1�΋� (u��q��������T1SVGUNYSɀo�'������ASK_OPTICONn�΅�������BCCFG ��΋O���I�2��` ;A�I�r]o�� �����8J 5nY�}��� ��/�4//X/C/ |/g/�/�/���,�/ �/ ??�/�/H?3?l? W?�?��?��0�?�? �?O�?&OOJO8OZO \OnO�O�O�O�O�O�O _�O _F_4_j_X_�_ |_�_�_�_�_�_o�X �  o2oPoboto�_�o �o�o�o�o�o�o :(^L�p�� ��� ��$��H� 6�X�~�l�����Ə�� �؏�����D�2�h� o������ԟR��� ��.��R�d�v�D� ���������Я��� �<�*�`�N���r��� ����޿̿��&�� J�8�Z�\�nϤϒ��� ~������"�4߲�X� F�hߎ�|߲����ߤ� ������B�0�R�T� f����������� ���>�,�b�P���t� ������������( ��@Rp��� ����$6 ZH~l���� ��� //D/2/h/ V/x/�/�/�/�/�/�/ 
?�/??.?d?R?�? >�?�?�?�?�?r?O O(ONO<OrO�O�OdO �O�O�O�O_�O__ &_\_J_�_n_�_�_�_ �_�_�_�_"ooFo4o joXozo|o�o�o�o�o �? 0BT�ox f������� ��>�,�b�P�r�t� ��������Ώ��(� �8�^�L���p����� ʟ��ڟܟ�$��H� �o`�r�������2�د�Ư����2��P���$TBCSG_G�RP 2���  �P�� 
 ?�   {���w�����տ��ѿ@���/�A�T�[��b��d0 �p�?�P�	 HBHA�L��͌�@�B   �C���϶ˀ��ϟ�D����A���x����A��T$�9��6f)f��f�@P�C�ώ�c@�f߬��C��� �߮ߴޥ���%��%� D�W�"�4���j�|�x������?Y������	V3.0�0s�	lr2c��	*2�*�O�A�\ ��ѳ33P�d���� x�J�y�  �������T�JCFoG ��l�Y o�����������=K
 %�Kq\���� ����7"[ Fj����� ��!//E/0/i/T/ f/�/�/�/�/�/�/s� ��??(?�/[?F?k? �?|?�?�?�?�?�?O !O3O�?WOBO{OfO�O �OP�<��O��O�O�O 0__T_B_x_f_�_�_ �_�_�_�_�_oo>o ,oNoPobo�o�o�o�o �o�o�o:(^ L������h�  ��$��H�6�l�Z� |�����Ə��֏؏�  ��D�V�h�z�4��� ����ҟԟ��
� @�.�d�R���v����� ���Я���*��:� <�N���r�����̿�� �޿ �&��>�P�b� ϒπϢϤ϶����� ���4�F�X�j�(ߎ� |߲ߠ���������� �B�0�f�T��x�� ����������,�� P�>�t�b��������� ������&(: p^����t�� ���6$ZH~ l������� /2/ /V/D/z/�/�/ �/j/�/�/�/�/?.? ?R?@?v?d?�?�?�? �?�?�?�?OO<O*O `ONOpO�O�O�O�O�O �O_�O__&_\_� t_�_�_B_�_�_�_�_ �_"ooFo4ojo|o�o �o^o�o�o�o�o�o 0B�oxf�� �������>� ,�b�P���t������� ��Ώ��(��L�:� \���p�����ʟ���  ��_�*��_�l�Z� ��~�����į�د�  �2���h�V���z� ��¿Կ濠�
���� �.�d�Rψ�vϬϚ� �Ͼ������*��N� <�r�`߂߄ߖ��ߺ� ������8�&�H�n� \���>�����x�� ����4�"�X�F�|�j� ��������������
 Tfx�D� ����� P>tb���� ���//:/(/^/ L/n/p/�/�/�/�/�/  ?�/$?6?��N?`?r? ?�?�?�?�?�?�?�?  OODOVOhOzO8O�O��O�O�O�O�N  PS V$_R��$TBJOP_�GRP 2��E��  �?�W<RCS�J\=��@0WP�Ry@T�P � ��T��T �Q[R	� �BL  �UCр D*W[Q�_��_?fffe:�lB �P�ff�@`�33D  $a�U3o>g�_�_�po�l�P�e9<�b>bY��?٪``�$o�oUA��gD�`$�co�Quz�9�P�Aa�P@>a���C�Z`Ep<�o]A6ffpu`asD/�U�h�͔r ��~�a�RieAq�`�q���@9q�|�d&p`%���c333D��\P8���?�`?1L�pAp[QB�b�k��}� ��z�� >�sffԁL���T� f��fo ��Nw@�*� 8�f���r�,���П�� ȟ��'����F�`�J��X�����SC�V�ء��	V3.0}0�Slr2c�T�*��TQ��� E���E��A E��E���3E�iNE��!hE�فE����E�I�E���E���E��rF�F��FM(F��5FBF�aOF�\F"�f,�z  E��@ E�� E��� E�  E������ E������ EȆ�Ԏ������ F   �F� F$ �Fj` F�@ �F�P F�` �9�IR9�o���L�_ ��V��LQ�8TESTPARS��XUP9SHRk�AB_LE 1�J[4�SV�+� �0�VǅV�V�WQV�	�V�
V�Vȥ�Q�V�V�V�뱅�RDI��TQ�϶���������f�On߀ۊ� �߮����ކ�Sl�RS 0ړ��������� ���#�5�G�Y�k�}� ������������/]k� o��*	�%�7�I��π��+�=�O؆�N�UM  �E*TQ�PP �����_CFG �����Q@<PIMEBF_TTq��RS~�;VER�<Q�;R 1�J[
' 8�RP� �@5  ��� ���//&/8/J/ \/n/�/�/�/�/�/�/ #?�/?Y?4?F?\?j?�|?{_�h@R
�<PMI_CHAN�G R �3DBGLVQ`IR;Q�0�ETHERAD �?�E;@�S ��?�?TO6V�0ROUmTe!JZ!�D��OwLSNMASK�0HRSAA255.��E��O�O8TOOL�OFS_DIq���5IORQCTRL �s[���n]8]_�_�_�_�_�_�_ �_o"o4oFo�
�_To�fo�og�PE_DE�TAIH3ZPON?_SVOFF)_�c�P_MON ��"P2�iSTRT�CHK �J^�mO�bVTCOMP�AT�h;C�d�`FP�ROG %JZ%�j�=?qqISP�LAYr��j_IN�ST_M�@ �|��g�tUSe]orL�CK��{QUIC�KME�0)�orSC�REF�3Jtps��or�a�f���2w�_{���ZyIS�R_GRP 1ξJY ؛  6�����;�)�_�M��8����Y�� �����͕�����/� �S�A�w�e������� ѯ�������=�+��M�s�	1234�5678����f�X�`�1�Ћ
 �}�ipnl/۰g?en.htm������0�B�X�P�anel setupF�}<�ϘϪ������� u�k�� *�<�N�`�r��ϖ�� ����������ߝ� J�\�n�����I� ?������"�4�F��� j�������������� _�q�0BTfx ������ �>�bt����3�~UALR�M�pG ?J[
  �*/!/R/ E/v/i/�/�/�/�/�/��/�/??<?�SEoV  �n6��ECFG ���m�6��A�1   ;Bȩt
 =?�s 3E�?�?�?OO+O=O�OOaOsO�O�Gz1ʂ҆�k SΟ�OH7I2sv?}{�`(%0?"_ p_I_4_m_X_�_|_ �_�_�_�_�_o�_3o��L� �M�OAoIm_E�HI�p1��i�  (p ���(/SOFT�PART/GEN�LINK?cur�rent=men�upage,153,1}o�o&3�'�o�n71�oq����6q);�eedit�bT��`�	��-� �)oS�e� w�������<�я��� ��+���O�a�s��� ����8�J�ߟ��� '�9�ȟ]�o���������è�R��aR��� �%�7�I�L�m���� ����ǿV�����!� 3�E�Կ�{ύϟϱ� ����d�����/�A� S���w߉ߛ߭߿��� `�r���+�=�O�a� �߅��������ʯ ܯ�'�9�K�]�o�r� ������������|� #5GYk}� ������1 CUgy��� ���	/�-/?/Q/ c/u/�//�/�/�/�/ �/?���;?M?_?q? �?�?�/�?�?�?�?O O�?7OIO[OmOO�O �O2O�O�O�O�O_!_ �OE_W_i_{_�_�_._ �_�_�_�_oo/o�_ Soeowo�o�o�o<o�o �o�o+?(?a s�����o�� ��'�9���o��� ������ɏX����� #�5�G�֏k�}����� ��şT�f�����1� C�U��y��������� ӯb���	��-�?�Q��<��$UI_P�ANEDATA �1�������  	��}/frh/c�gtp/whol�edev.stm�c���ӿ����)Gpri��.�Ip}2��V�h�zόϞϰ� ) ���Ͻ������0�� T�;�xߊ�q߮ߕ���p�����Bv�Nq*�=�B�T�f�x�� ������3������� ,�>�P���t�[���� ����������(�L3p�i��  ��������� 1C�g���� ���L	///?/ &/c/u/\/�/�/�/�/ �/�/�/?�/;?M?� ��?�?�?�?�?�?0? Ot%O7OIO[OmOO �O�?�O�O�O�O�O_ �O3__W_i_P_�_t_ �_�_�_�_Z?l?o/o AoSoeowo�_�o�o O �o�o�o+�oO 6s�l���� ���'�9� �]�D� ���_o�oɏۏ��� �#�v�G��ok�}��� ����ş,������ �C�U�<�y�`����� ��ӯ����ޯ�-��� ��c�u���������� �T���)�;�M�_� q�ؿ��|ϹϠ����� �����7�I�0�m�T� �ߣߊ���:�L���� !�3�E�W��{�� � �����������r�/� �S�e�L���p����� ������ =$a����}�r�����)�*�� Vhz��� �����.//R/ 9/v/�/o/�/�/�/�/��/?�������$U�I_PANELI�NK 1����  � � ��}1234567890_? q?�?�?�?�?�4��]? �?�?OO1OCO�?gO�yO�O�O�O�OYIY0�:�M��[0-/S�OFTPART/�GENA1?CON�FIG=SING�LE&PRIM=�mainedit �OI_[_m_YJ_$_�M=wintpe�,1@_�_�_�_XK  �_$o6oHoZoloo o�o�o�o�o�o�o�o 
2DVhz� �������.� @�R�d�v��� ������Џ����M 0�,M9P E=Po�r?S�,Ico :�{�^�������˟ݟ �����7��[�m�P������O���BS0ߢ��C���/�%� 7�I�[�m�`C����� ��Ϳ߿񿀿�'�9� K�]�o��L���э͙� Q|����������!� ��;�M�_�q߃ߕߧ� 6���������%�� I�[�m����2��� �������!�3���W� i�{�������@����� ��/��Sew ����.���z� !E(W{^ ������/� //A/���͡Ϸ�}��� �/�/�/�/�/?�2? D?V?h?z?�??�?�? �?�?�?
OO�ϝϯ� dOvO�O�O�O�OE�O �O__*_<_N_�Or_ �_�_�_�_�_[_�_o o&o8oJo�_no�o�o �o�o�o�oio�o" 4FX�o|��� ��e���0�B� T�f����/������ ���ُ���>�P�3� t���i�����Ο��O/ �s/(��/L�^�p��� �������?ܯ� �� $�6�ůZ�l�~����� ��#O5OGO�� �2� D�V�h���Ϟϰ��� ����u�
��.�@�R� d�v�ߚ߬߾����� �߃��*�<�N�`�r� ����������� ��&�8�J�\�n���� ������������m�" 4ßXjM�q� �����B T7x������ A��//,/>/P/C� t/�/�/�/�/�/�/o/ ??(?:?L?^?Ϳ߿ �?�?�?�?�? OO �?6OHOZOlO~O�OO �O�O�O�O�O_�O2_ D_V_h_z_�_�_-_�_ �_�_�_
oo�_@oRo dovo�o�o)o�o�o�o �o*�oN`r �����m� �&�8��\�n�Q��� u���ȏ������"���?�?�{��$U�I_POSTYP�E  �5/� 	k�{���_QUICKMEN  ��j������RESTORE �1ו5  ��/
�2�D�h�mc�������¯ ԯw���
��.�@�� d�v�������W���˿ ݿO��*�<�N�`�� �ϖϨϺ����ρ�� �&�8�J���W�i�{� �϶��������ߡ�"� 4�F�X�j����� ����ߋ����y�+� T�f�x�����?����� ������,>Pb t������ (�L^p� ��I��� //ވ�SCREܐ?��u1sc�-�u2M$3M$4�M$5M$6M$7M$8<M!��USER/ 4/2F"T. O#ksW#�$U4�$5�$6�$7�$�8�!��NDO_C�FG ؜�  �,� ��PDAT�E �)��None V��S�EUFRAME � 
��&,1RTOL_ABRT7?���N3ENBX?I8G�RP 1�!��?Cz  A��3�1���?�?�?�?�?FO"OG:ېUx81g;?MSK  {5�A�g;N41%a��B%���O��VISCA�ND_MAXyE�I�c8�@FAILO_IMGy@f����#�8�@IMREG�NUMyG
�KRS�IZyC,���$�,SONTMOU4W0{D�%�VU�#_�c�� �P�2�FR:\�O �� MC:�\XS\LOG�VB@4 !�O�_�Q��_o
�z �MCV�_�SUDM10fEX9k
�f�TwV�2ۜ��p(��o=��͓o��j �o�o�o�o�o�o�o  2DVhz��K_PO64_?S�0Π�n6�uQ0LI� Q�z�x�qV� �|�f@�w�� =	��xSZV�~�����wWAI��DST�AT ܛ;�@�_ď֏�$����E�P12DWP  ��P G/����q��AP-��B_JMP�ERR 1ݜ�
�  � 2345678901����� ��ʟ��ϟ��$�� H�;�l�_�q����LT@MLOW���P�@�Pg_TI_X�('�@�MPHASE  �53��CSH�IFTUB1~k
 <���Ob��A� g���w���ֿ����� ����T�+�=ϊ�a� s��ϗϩ�������π>��'�t�K�!��#���:	VSFT1֣sV�@M�� ��5��4 �0��UA_�  B8����E��0p�����Ҫ�ӌe@��ME*�{D�'����q��&%�!�M��$�~k��9@�$�~�TDINENDcXdHz�Ox@[O��aZ®�S����yE����G����2�����������REL�E�y?w�^_pVz�_ACTIV���H��0A ��K��B�#&��RD�p��
1Y?BOX ��-�V���2�D��190.0.�� 83��254��2�p��&��r�obot�ԟ   pN g�pc� �{��v�x���$%ZA+BC�3�=,{� 낆;-!/^/E/W/i/ {/�/�/�/�/�/?�/ 6??/?l?!ZAT����