��  L��A��*SYST�EM*��V7.7�0107 10�/3/2018 A]  �����ABSPOS�_GRP_T �   $PA�RAM  �  �ALRM_RECOV1�   $AL]MOENB��]�ONiI M_IF�1 D $ENABLE k �LAST_^  �d�U�K}M�AX� $LDE�BUG@  
�GPCOUPLE�D1 $[PP�_PROCES0� � �1��U�REQ1 � �$SOFT; T�_ID�TOTAoL_EQ� $�,NO/PS_SPI_INDE���$DX�SCR�EEN_NAME� �SIG�Nj��&PK�_FI� 	$�THKY�PAN�E7  	$D�UMMY12� ��3�4�GRG�_STR1 � $TIT�$I��1&�$P�$�$5&6&U7&8&9'0'�'�%!'�%5'1B?'1I' &]'2h"�GSBN_CFG�1  8 $�CNV_JNT_�* �DATA_C�MNT�!$FL�AGSL*CHE�CK��AT_C�ELLSETUP�  P� HO�ME_IO� }%:3MACROF2�REPRO8�DR�UNCD�i2SM�p5H UTOBAC�KU0 ��	DEVIC#T�Ih�$DFD��ST�0B 3$�INTERVAL��DISP_UNsIT��0_DO�6�ERR�9FR_F�a�INGRE5S�!Y0Q_�3t4�C_WA�4�12JO�FF_� N�3DEL_HLOG�2�jA��2?�1k@�?� ��� �M�OTOR_CE 	 h Y0M_C� � �	�BREV�DBI�L�GGXI0�BR� 
 [ OD�<0�A	$NO�� Ms0�@�DR�!�YW �VAQ��A_D�# d� $CARD_�E�@T�$FS?SB_TYPi� �CHKBD_SE��5AGN G� �$SLOT_NUMZ�QP�A�C��G �1_EDIT�1 � h1G�=H0S?@f%$�EPY$OP�c iAP_OK�sRUS�P_CR�rQ$�4�VAZ0LACIwY1Db�P|k �1COMMEc@$D@fVa`�� ���QL*OU�R ,�@�1V$1AB0~ OL�e<Pz CAM_;1� xCQg$A�TTR��P0AN�N�P�IMG_H�EIGHrQsWI7DTH�VTCRe��0F_ASPE�CrQ$M@EX�P;$� Fv�C�F\T X $�GR� � S!1NpB_@NFLI<pwt
�UIREs3��QO}MqWITCHvsJQpN.0SXt�cG0� � 
$WARNM'@f��P� sLI? �qNST� �CORN��1FL{TR�uTRAT@0�T�pAP$ACC��1�  �� �OR�Id`|S�{RTq0_sSF� �!CHGI1RTspu3MII�TY�2p�K*
2 �`�p� 1sR*HD�cJ* �ȁU2Æ3Æ4Æ5ÆU6Æ7Æ8Æ9���*�CO�$ <� l~�x�s1��`OIT_ 2 w 4� STY�rw2Ge!VAR���)Y0���P��p��$ ��P��2�@�2�0D+P��0'`?�OJ�u4TOCO�3PE��USH_�CEp�p������EXT9��E�a�E� 1 2� 
��.� ə 2P����2@0>��  Hip� Q�@1𕃗�p�4O O���q_�s�0o�� A~�ʘ
:�bM<��r��g��@n�TRIGz�dP���@0��j@A��5�P�6������w�CO_MO�Rx� tW�FL�Ev�NG�1pTBA� .s㴴Q꺸�߸VP�BQ��P��0Ż��w�p�`�P�2� W�%��J�%�_R�k�hPr�J�(�vȑ�J��D�C����}�w�ul�P_�}0OF� �  @�� RO����PqIyT8C�NOM_�02�1"�q3"���$� �4����xP٥}E�RAG�0� �0��	�?R
$TF\����MD3�T��&@U=0��Pb�H,�2{�T1��E,�� �u��v��v���OPDBG4q� U��`PU�����4���:�AXc��rbETAI�3BUFnV��)���!  |�p9��pP�I�b�P��M���M��+���F��SIMQS���҂aP���!�8�Cµ!~���@~0JB�pL�}1D��A���@�-����"� � �PNS_wEMP��$G��Ą��P_��q3�1_3FP:���TC��9p �r��q0�s���ӎ�� �V�QAR�!h���JR�!0ARSEGFRA�'�v 0qR�T_LsIN�S$PVF�����,�#2R�D���a*)B��F�$( '�Ϝv�u�cӳ�a�=�.0m��M��	=�SCIZ$� ��T����

�aRSINFz����) �p��<
 <�� Lh��Ў��qCRC�uFCCC �pr
 ���}��Lr�A���q��]�D�t�s�C�j@֐��`$ pP�ٰ+(EV+&��zFA!_��F��N�m&����b����#A1���!% �.�s߻RGG`��)�F �b��D<�24�LEW �As}Ұ���.SP�`s&x 3�E������Q�R���`Ch�$LG �p���1Z`ѰlP�Pq!A?@ٰ.�Z�R�"����3P�s�3)�8RA���3AZ���8' �ՍOd�FC�bApQpF�p�4�)�s�ADI LKWqOE�0/r�0ٱ�p >D�p�p.s��S�Px�L0q�QMP.�`YCH��0���U�baU��]'��TIT�!�S⑕%V�n��DBOPXWO^��(���$SKdюR��D�BTf0TRL��)�˲A&`���0�`��DyJ�ā�_CAL�Q0bWPh@_WPLnLa�ߒD�a|W�a|W��!S�1��*R��PRc 
#P��v���g+ ����$��{$� �L�Y!,�_�S���-�_d�� .odENE��!/;o�S�P��ORb0H �b�On +$L�c,$�S���0�k+ 4��ձO�0_DwA��ROS�r��[�d�Z�d�cN�G��ePA+�|[�/ETURN�bv�MRt�ATU�pvB�CR:�EWM=��GNAL����$LA��Mu;�-{$Pj�.$P@F��/ap�Q�C|t-ӶDO7 j��d�a|��fGO_AW��Ƹ�MO�p�B��DCS��1<mQISZ0�@֣�@@���r5�qDᣐ�r@������q��qW���NTV���rVE�}���w�f�փ��J�m&�����SAFE�9ա�_SV�BEX�CLU�����"ONL��ȃY_�y��=En4HI_Vv@��PPLY_�m�VRFY_[S���rr@��_ 2a`P�ќw��� m��qS�Gz  3R�
$ $�*pGq�� X�;����B���V[�u�l�AN�NUN碓��ID��U�bŃTp� ��б�b@��Ֆ�"QEF��pI5b4�$F����D�OTJp�a� $DUMMY �Q��� �#Pm0��u5 ` �HE�6U��W�уRrk �SUFFI	���pZP�!nP"�5�6�=�"QMSW�u6 =8�KEYI�-�TM�a�ӡ,qΦI�N<�հ!Rr@�t7 �D��HOST�P!��P��� �����EM���k��P�SBL� UL�R8� S�6z�=�PT�|`Ʊ9 � $<���uSAMPZ � ���D��O I�`H�>L�$SUB�����4`�]ၲ�C��SAV������ �3s@�,܀��P$`E<AP�YN_B
S: 0&�DI��nPOU�F�v�C$��R_I;� �ENC2_	S�0P;Qs@����1�¸@Ń��-pBQ<R�����a��>��=  ��z����`pK�ddAn���AVERˡ���(��gDSP���PC8����B/�Uѣ���VA�LU�HE@�M�X�IP����OPP~0 .�TH���#��"}�SY@-Ս�F;���ad��w��@.SC8�����ET�$>���FULL_DU ����Dp����1g����OT�BM��`NOA�UTOQ?	�$�R�S���Q�CJ��a�C>R/0��O�L @H *a�L�@�#� ����$�`�������� �Q��<��校�櫡��U7��8��9��0����1��1��1�1��1�1)�16�1JC�2Q�2����2��U2�2�2�2)�U26�2C�3Q�3��3����3�3�3��3)�36�3C�4�Q�D0SE�RA� <11�'S��Â1I`��^�v��FDӐ��B L�V1�!�V2]� ig��-REG&�UFE8.p8pPC ,_���? �p�0?(�к�E�p�Т��"PD?�$�TPA$VARqIg��UP2*�3E 0���TD�����#x��,'&%����B;ACRF T�����D)�L���P� IFI��P� �@<0~%5P;Be`�F)p��>PGt ;���2�� ST���!�@a� �`�&�/0	�"C+4	7P���s1�%�1(� 47FO�RCEUPl���F�LUS�H�Bp�_�E�2�D_CM�pE��h45IN_pY3m�^�
8REM]FŁ71�5�P62�0�8��:K�9Nw��8EF1Fӿ4�pINC�62wOVMIOVAI�TROV<N17DT<�HDTMXkL�0 H�pkJ҆P�H�5�C,�P62CL0_���Jȱ`k��9_Q��8_T�k0�KQ��pAL�Dz@42 X���Q�6�F�Xa`RQ44^IT�_�-�#0M"E��C9L��ıRIV���nREAR�IO�5#PC���@7B�r
8cCMJp0� dA�GCLF+S�QDY��X�@ב�S5T�ED�G01"E`e-GS9S�P�H P�=a�a����_<aSh<a�1��E�c<a3uk5�uf�GRAE �$I� ���W�ON<��cBEBUGp��b��4��p��_E �J ��D ��TERM�eK�iO�RI�1�`L�f� S#M_ꀹ��`M�eI���TA,yN�e���UP��O� -��q��Ju��cspK�$SEGxz	`ELUSE�pNFI�!�r��a%�tot�L$UF}�H�!$U����p(�A�w�`T��� �NST��pPAT��a��PTHJ��&���V�r�5���up��J��qR�ELN�-�SHFT�Ңq�@�_SHOQR	�#�+v 6p$Ewr��N1� OVRjӤ-���Iq�qTU� �AYLO��RC��I�R[����h��ERV��݁0����w��pN�w� 8��� Rz�QPi�ASYMu��i�qWJ�w�&PE �<�h��)�U���p B�@�p�(�V�Ph���,hл�OR�pM�#L�_GRSMT�%P`�cGR5 �c�PA�p����� �Q � u�(r!TOC�q��P��� $OP@�"(���
� DQYOR1ӰRE_�R�sP-����� ef�R��z�X�x$e$PW�RZPIM���R_pU�{���r R�b�Hi% �_ADDR~H_LENG�P��
�M�R00SH�S HS��;�w�I��I���I��SE�[An��S3�#T� $��M�~1_OF�F[Ґ�PRMU� �'�TTPu_T�H��U (��OBJ�R�x$$�LE�ĳ��V� � ��AB%_!QT��S�q36� LV��KR�R���H���BG>�LO0��	Q��p�Q2w�̜'x�SS@��HW�=�q��WD���I�NCPU�bVISIO��-�����_����m���� �IOLUNZ"X�UPCb1�$SL���0P7UT_Z�$���P�P"���~0F_AuSCbY` $Lu �u!���0U+p���q`��e��߀HY0��fӢA�UOm0BcZ `RЫ��B}��@���ѧ�Pq3�����ф�������UJ��&[�!NE��JsOG�w,�DIS2b��K��	0Bc\ Q���qV�j�CTR<R�j�FLAG�bG;LGAd] �0P��ҶcLG_SIZ��5 �� ��I���FD��I�������  p���q���9�� 9��I�9���9� p9�z@S�CH_/ �Ŋ��L�NK��^��v1E Rb!��� U����r�L���DAU���EA����A�����GqHB���U�BOOZ"�_h Al�� I�T+�`h�REC�1
SCR�0<�m�DeIg�S�p00RG�" �Qh5�`�`��W�U�	S��T�WoU���`��JGM�MNCH|�#U�FNKEY��K�PRG�	UF�����FWD�H]L3STP�
V���p�# �RSkHԐ]�C��I��`��P��U���������u�G�	i�P�O'N^IM�F�OCU(RGEX.\�TUI�I�{"��#��#� ���A�P�R�N��O�1�$ANAUқrsPoVAIL�CL�Q~l�DCS_HI�d�2_�2O8�Q4S�=P/58S+8�IGAN�� �����Ta�N_BU@@�`e�5ĀT�"$��FP����r�s��2g�ae�Ā��ü��p" U1�52�53�1'p�7"0@�b � �����u(�B(�ID$_@�P؂��O@C��qNFST��R��Y�&p��q@ a$EFCK����F�F8��7$c L��{� �`�؎�X�g����j��駨O_ d ���c�O0S��`C��e �@C�LDP��l�TRQ�LI ��:�dYRTF�LGzBRP�a�S�!DY�W��LD�UpT�UORG:��R�����X_��m�BT�df A��`pT�aT�US�	TdP�``�P?dja>JcRCLMCUd�_��_gi��Ga*�M9It��g d��"A�RQ�c$DSTB�:�E@ �f�hA�Xl� �h�lEXGCES�r���bM��
hP�bl�v��j@�i���f_A�j���X{�o�hBPK��j{ \��GROU��n��$MB��LIܱ~�sREQUIR�r�o��|O�{DEBUT"qL�@M\�k
��m����sUbqND��,�@�l���o�fB�DCI"��INʰ@������L�\�W0N8b�q���`@/�PS�TD� m��LOC%FRI��%E��%E�A"�&A�aqODA�Q\�n X��ON��F����	�KI�B�U�U/������AFX�`IGG/ o �`�Cq�<��C��DR0�%oCk����{��Њ�wpu�DAT	A�7ǐE����q����N�2p t $+MD�Iݱ)��C0��a��H؀$� ��<���ANSW`��(g�W!�D��)���=`@�q +pCU���V?��P��RR2��r Dհ�.�A�Da d$CALII�`R�G�!��2���RIN��<��NTE
��2sy��8�X���
�_Nt�@����a��Dru�7DIV'�DHp�:ve�$V��[�vEA$�$Zӂ��Q�0ӂ�����w�H �$BEL�Tn��AACCEL�C1����ŰIRC��Ѐ�Ф�TcA���$PSpWRL�0 }���lS�۷��� ܶPATH��1�ѳ1�3 �q_�1��b��h�Bb�0C���_M=G�$DD��ܰ_$FW��ڐ�����ѳ����DE��P�PABN�ROTSPEEx��1��"`�J���1D��`���0�$USE_���#P����SY����Ba �r�YN�`A O�OsFF�O�MOU��3NG�"�OL!�|�INC^�Ձ�¥��bx�׀`�bENCS������b�����d��IN�WBI ���@�Gb�V�E�Ы��23_UyPy��LOWL71A�C�"`��3�D�@�b�p� P��erC�����MOSd0|tMO���/pBgPERCH  P�OVG�KҒ� %A��pA6�EdpAۃ�� �`�p;�?�40Ve�Wp���L�$��yw�����UP����1�L�TR�K��SBAYLOA 1Q��Tqa� �p�e�րd@��RTIXq��d@MO�����bTr�P~��d�ç�|�3��2���DUM2\�S_BCKLSH_C � ��r�q��WӉ����
fѨ�HaCLAL��0��+a��#@NCH�K"`[ESx�RTY@L�#�ӭ5�Qّ_jCNf�_UMXp�	C�Γ�SCL���LM?T_J1_L�P�`�(��E�� �p� ���SPC0k���9��PC����!HP�p�šCc`RsXT����CN_¢N���ѳSx0F���V9�ZC�շ�m ��2qC�0�SHjC¢ �����Q���֣�d���>%���PA���_	P���_eP� h���0"ax�${JGw2}$�!�OG���TORQU+�ON^����`�r|������"_W��a�_q�5w�5}�5UI;I#;I}�F�� 1J�ab8a��VC"��0�d�b�21�>p8�?�b�5JRK�<�2��6=`DBL_SMt��;bMY�_DLw�;bGRV4Dw�D}��1H_P#�34�;J�COSHK��HHLN �0kK�5rDw�mI}�mI ?1�J�L]1�5Zf@|���1MYtA�HTBTH|ZMYTHET0<�NK23}�2Rq�u@[CB7VCBq�C�a�r\R?4jQw�jQ7VSqBw��RBUGTS4q��C�!Ձ?#�DV �Tx�C�W�C$DUx  yx�Q�����b�V���a9Q��ۆ$NE1t@�AIv@��U$�$U�&QA*USe\g:EEHEA�LPHXu1b�1bS �5�c�E�c�E1b�F�c(�j�FU�VuhVjhg���lV�jV�kV�kV��kV�kV�kV�iH�uh�f�r�m!�x�kH��kH�kH�kH�kH*�iOflOuhO ��nUO�jO�kO�kO�kUO�kO�kO�FF1b�WQ���E��hgSPBALANCE_�A��LE�PH_*US�P롈F��F��FPFULC�6��6��E��1s��UTOy_s �%T1T2w���2NZ�����&�@��8�`²���T"��OK�ı� INSE9G��U�REV��U����DIFK��1tl�I�1u �OB��>CǩMI�e�4?LCHWAR�²��ABZ!��$ME�CH`Q�@�t��AXn�P��LgX�l��v 
���!����ROB��CR��Х�;��SK_�_x P ��_)�AR��x���M�1�������V�I�Nݑ�MTCO�M_Ct0��y � ��
���$N'ORE��i��F�X�7z 8� GR�"y��SD(`ABz�$?XYZ_DAia���DEBUݑ}�F����{ �$G�COD- Բ��z����$BUFIwNDX�  ıwMOR��| $a��Uɱ]���v���7�G��} � $SIMUL� �۰���T���OBJ�E�T�ADJUS<r�e�AY_I�!���D�ǻ��w�_FIz�=�T� ��� �ǯ�*��������p:��DD�FRI���MT
RO� ��E1z-��OPWO�0���~0�SYS�BU�`��$SOP�L��SW�UV��PgRUNH�}�PA��D|�x�Q���_OUb�1q�*���$��/IMAG-��`�P�IM/���IN��0����RGOVR!D��n�]���P�����)`L_j�� ���RB�*`2ML!?�ED�z� "�NC�M^�!6���S�L��� x �$OVSL��SDI*�DEX�����m1����V0��N ���!������������M!A)u�_SE9T� ��� @� �L��RIV��
�!_dQ �9�,���|p�� � H���y�z ATUS��$TRC`����t�BTM}�g�I�����4 S�\���� �D��E�Л�q�LpE��r��: > r�EXEx��D������	�1�� �w�UP����s$+���XNN���m1��|1�� �PGnV���1UBf��6�f�:�JMPW�AI�P��~LO�� a�F�S�$R�CVFAIL_C�aЁR������}�� �Ű��@R_P=L:�DBTB�!��a�BWD�q�UM� �IG���Н� GTNL�� R�^�E��H���Q �DEFSP�� G� L����g_jx�xUNI�Ӣ�vb#R����@_L�-Pp��PI����а� v����ర��:�N'�KET�����P��� h~��ARSIZEؠМ ����!Sp�OR~:�FORMATc��
COz�!ߒEM2��4$�UX;����6�PLI��� � $S�P_S�WIG����0� A�L_ ��uAR-�BB�\PC-�D�ѷ$E���� C�_9� � �c (5-��!J3�P�-�+�TIA4�)5:�)6-�MOM)�	3�)33)3#3S�B� A�D	3M63M6#3PUkPNR.4z53z5#2�P�x"���� A$PI(f�%��$D �5!C�5.C�5mT�6�; �T�T��V��ܡ��|��SPEED�pG�"ZD�gaFg� � ��aF�CpH�I��SAM����DaG�C�MOV��TQ@���UTeQg1;�/T2;�%�*�0U� 2��H��SINb\�  �CiX�[`T�kZ�X�T<�[�[GAMM߆a>��$GET�����|�D�$0�
��LI�BR7I��$H�I _�р��@fEĲ MhAGnj`[fLW Bm�flji�f[f�"���H��A� $�PDCK;���|�_�@'�0�^R�)�!QU�w)3tM6y�# ��$I8�R��D`.�V�!�X�LE8�`�@�x�(Yp��u%�4��0�PґUR_SCR)�q��C��S_SAVE_DX%��uNO� C@� �$�pd�*�6�O� �9���H�8���.�'F u�EP�!���@b�U 8W$R<�[HQ�kF�H@هՅ��Qt$M�5� �!�QW���@2s*����p���W
�آT�J�`�~0H�r2�MŰx�CLw�w �M�qC � �$PY� @�$W��[�NG���!���$ ���$���$���$� +à=�#`�#|�� X�O��#�!Z+�w ����# p��S�3s�6�@/�A�S�e�@��!_Y�� |���)�p)9� 3�#3�p:���:AE��e��ä�r����� ŤP$!�PM���QU�@ � =8�QCOU5qa�wQTHƠHOL��oQHYS; ESQF��UEw��r�OT�  �Pd�8e@�sUNy�z� O 9O�°0� P��ִp��q��7ROG?���;�2��O �յ�ü#���INFO?ѕC ư�I�:�ȿ�OIL (KpSLEQRFt�FEt��$��D� �0����`QO�`PSC?aE}`sNU�Ǿ�AUT�q��COPYQ �����M��N������C��>� �RGA+DJ��"XS��C$�W�8�W�WU؁PU؍pW�jCG�kE�X� YCӒ�R�GNSS� ��$ALGO�c��NY�Q_FREQ��W`�PEF��I$>�LAus���S�$3�PSECRE� ��A�IF���NmA�A%&�_Gusk�Q�˸Tf� ���*�R��P��mr�4���ELEr  � ���!NABӒ� EASI��قRN���@SA�q��NP*`I-��t��iq��� �s�AIBx� E�n@VXp-�BAS�"/�*bu�TR�� �Q��$F�n�c�c��ip��~�� X �� 2��U�T��x����w������$�2MPO�W�M ǰ_B�!��
�	)�>�ԝ � &�� p��3�64SRVF�1)S��C T_Om �\�3�	��5*�	6�	7�	8k�ѹS�r�0� @�M�C_F��<!��L�q�q�Y�R��� hP��3P���� ,KpFLА�q�pSYN� MM��C��PWRU�P��0=�ĲDELA�F�Y� AD���QSwKIP�5� �C װO��NT'Q��P_װ ���p��� �.C�;C�� ��  �� �� �� �� z�9hq�J2R^@n�0� 4��EX`T�ӎ!=�ˁ�!��Rp�!'�R��RDC��ף ���R_�OR�v�FUpQ�*���"�TR�GEAR�亃mrFcLGl��ƠERr��C<ç�UM_� ~{�J2TH2N�3~" 1� �!uG��T�` �R�w0M^1]�I�D�REFQ1�q� �lQ��1��_1ΐTPEbp��EG���� �1��S�2ݳNb5��2�О42�2��?�?�?P�?�?OG3�2�)O@;OMO_OqO�OG4�2��O�O�O�O�O _G5�2�#_5_G_Y_k_}_G6�2��_�_�_P�_�_�_G7�2�o@/oAoSoeowoG8�2��o�o�o�o�o�oESSMu�̠�n03�ʟ3E�q\��0MOO༴�� ��r��Lˁ�sIO.��yIUp|ˀ�sPOWER�� _�L�!��Ơ�̠�G�$DSaB��A�9�W�RTzyC^0�uS232�u����T�DEVIC�EUH�̈́ʂPAR�IT��W�OPBI�T����CONT�Rްˁ�1��ʂCU����UXs�s��0ERFACr�Z�[���*J�CH�Ѳ� L������C�>�EFROM��{�GET_� k������pTu�ȔJ�P|Ӏ�ѳ� !x$USAP|�(y��Ы�4�O���R�8႒,�_ONP8{�����WRK;M|��ὗ��SvFRIE�NDF���$UFx�����TOOL��MY��$LEN�GTH_VT�FCIR��+���~�E@��9�UFINV*� ;�qRGI��v�OAITI�2�X�lA���G2��G1�0~�����P�����O_p�������$�C��	�TC?�A�ȡ�� �G*0Z��д� s�p�󪞘W��W�Ѧ�p��E��OX ]���L��T��H( ���О�p�$C�R�W������ɴD���`���ٱL��$���pH���0��1ʘ��2��2-�3��3ʚ�t� ˙;ɐ�Sv��\���h�S$V� @�V��V� (���ж� چ� �pb󦲂 ����c���V���V�?��1au3$A� D�PR� E�D[���S!v�)!�B��ҷ 0Io����� �ķ�pC��ԏ0�
��S�q�� ���RY�����$RUNN�pAX���A�L&����/THIC��K�|:��1FEREN��>��IF_CH����aI��E�Sv��G1`��d�Rpk�����_J�F��PR����RV|�A��2}�2] �VAL�  ���� ��r��  2� �S� ~U��d �$E0z�5L2GROU�q��TOT���DSP,�JOG�񖂷 _P���O�� �A�ĆK4�_MIRȗ�j�ȠM����AP���`EP0���M1ScYS�s�M1PG���BRK��,�,�Icqp��������ADՁ��BSO�C ��pNDUM�MY14����SV���DE_OP��S�FSPD_OVR�/�C� WZ�OIRe5pNk�fF,�lfE�OVH�SF�
�О^�F�t�l�̣8��s�LCH}�RECOVV��E��W�ME H�ROȰ�(T�_���� 9@22s�VER����OFSs�C��w�WD	{(h���B �TR���q��E_�FDO��MB_CiM�q�B8�BL��h���r�V ���&��-В3�G���AM������0/_M����)0�s=8$C�A;�)0D��B HcBK*��W!IO��qf%�q�PPAZ*��!k)�$~%%�r=DVC_DBv��!:� %�� t��%1�*0#��%3�&6ATIOs��2s�VU��:��vCABQ�ѣ���G��E�_���S�UBCPU$�R�S Ր���+�\��7���� ���$HW_AC#@����7�A��~��l$UNIT��}l�1ATTRI<���2R�CYCL�N�ECA,2��FLT?R_2_FI]�9�23+�LP^�=�<�o_SCT��F_�7cF_�<BJFS*���2CHAՑgG�A8����BRSD:&��	�%��p_T�PcRO0���EMkp�_%��8�B�� 1�B��3UDI`��?RAILAC�#7�M��LO �4���(�661�650#PRJ� S��ОQC�!ze�	/FUNC��>�RIN%�-���HP̾T��RA�PA� �B �S�P$�SWAR�|�C BL ��WdA0kAhhDA���QRhceLD�J ��zc���Q(�zcTI�0Қe���$v�R�IA��t�AF�0P|��c(�e:�߲�#�NCMOI�0�DFa_$��'��LM�{FA�HRDY��ORG`H�@����|Z`uMULSE$�x �7�� ���RT���p$�m$��$� ��|��U��� x���EGG��J �qAR'�;3209���u>`���AXE/�ROB�,�W~���_�}S�Y���q���S$�W�RI��|1;�0SCTR+�����q E�1A��M�zS����Bq�`<x���2  OT}���P	$(ARY�,�hQ4��]�FI���s�$LINK(q�ρ��_n�<�L�y���XYZpZ! ����OFFDR΂�����B*���RT�P�PU�FI@n���MB�TE�_JW���oۃ�O�P_����5����T�B��WrݒCB@��D�UZK�6{UTURN��0�����Q��H"ŗFL��� K3�p4���t�7<R 1����KQ�M�K�8�{U�50Қ7lORQ V�Q�Sv��s)���x�
p1��Us7�T��OVE ��Ms@w�}s ��s��r�W�M1 ��0���PsA�`� ���Y��"w����`���s��>��QERV�
�Q	REA���S�A����r��UR��YaV6YaAX��Ya5� ��9���9���9ǀ�F� ֐F��F�n�Fʔ�F� �pF�S�F�pC�pS� pc�ps�p��p�� p��p��p������oDEBU�3$�Q �a1T��Y򂏗�P�PABYWW!����HP��
���#��մ1�� ���-���֑����� n��ה����q�d���b\ЂU�LABk�ť��0�#�:�  ��pERVENB� O� $0��PA�!��POKO �x�����_MRA �� d ��Ee��ERRC;C�`TY�@%�IJ Vk�5��'TOQ4�r�L�p5��@����0C�q � p��T����E0_V1��7�_�;Sl�2e�2t���x��8����~#$W$@��j?�V�q���$�@R�`5���?�Z	�pFZN_CFG�p� 4�0w��@���3'�x� �` �����s� � ���@	$2q���@`�FA�`���fdXE�D�`	/��q���0�PM2�pHEL�L��� 5�n0B_BASY3R�SR���P�sS��1�a� 1��%�2�3456�78�ROaO�`Հ��NL�q��AB��QP� AC-K��IN��Tr@i1�萾�Pp�A�_PUfYCCO�p��OU��P
`
aP�@BU7�TPFWD_KA1R�� ��RE��/pqP0`a�`QUE��P�B@L4CSTOPI_AL������^S��3����SEMȤ3�$�3M�@� TYf�SO� TtDI��
@"`!U7�a_TM>�3MANRQ�&���Ec@Ss$KEY?SWITCH^SAA��!L4HEB@BEAiT"Q�QE�pLE
�TI8U#F�$"T@�%�O_HOM�`On�SREF�PR�QP&��^��Cc0OyC�`ECO�ි�`�`�IOCM�p'�!����p@��� DH��2 U��^"M�bx4"��FORC#nc "�7OM�p � @���c�@Ud�P�p1eF�T�p�3eF4��NPX_�AS�� 0 A�DD2 4$SI}Z!$VAR.MpTIP��Cj@AKB���S���@�2$�P�rS"�qC�VOFRIF%���SH ZI�4�@NF�"�p� n��� x��SI#��TEO�Ԣn�SGL`QT݂@�&$0yS��<,�aPSTMTM��S�P�pD�BW�bTS�HOW�U&��SV|p�t�� ���A00,�ٱ�Rn@�W@x@�W�@�W�@�W5�YU6�Y7�Y8�Y9�YA�Y�p�WY@�W_��V{��WF�XS��h�Y�� �hi,��h)i��hCi����h]i1ji1wi1��i1�i1�i1�i2��Y2�Y2i2i2�i2)i26i2Ci2�Pi2]i2ji2wi2��i2�i2�i2�i3��y3�Y3i3i3�i3)i36i3Ci3�Pi3]i3ji3wi3��i3�i3�i3�i4��y4�Y4i4i4�i4)i46i4Ci4�Pi4]i4ji4wi4��i4�i4�i4�i5��y5�Y5i5i5�i5)i56i5Ci5�Pi5]i5ji5wi5��i5�i5�i5�i6��y6�Y6i6i6�i6)i66i6Ci6�Pi6]i6ji6wi6��i6�i6�i6�i7��y7�Y7i7i7�i7)i76i7Ci7�Pi7]i7ji7wi7*d�7�i7~�7�d�2�VPG0UPD���  @�0���YSLO�� � �E� ��4W�G}0�հv0����ALU���&CU����F���ID_L�#��H�I��I9B$FILcE_�"�$$�3v��SA��� h��~N�E_BLCKK#�[�{Qd�D_CPU tٳ@t٧@%�7Ԃ¼T0�R �P�
�PWOP� ��L�A/2S��������RUN~�������0�~�"���"��� �T�BC�CE�Xw -$I�LEN�# V�#I����I�! LOW_AXIK#SF1I��2��M����|BP�I� ,��TORQ!I���D���?PLu �2��pI���[0_MA�@p������TCV�>���T�!?�^�T� ���������J����M��� J'�P������U�2�/0�������q JK��VKС!�!3��J0l
JJJJAAL
@ @ :e4V5|^�N1e�Pq 0���L��_�Q��P�1E��� `X�GROU��|Q�"}BG@NFLIC�C�� REQUIRE�4EBUy3E���@D�2��AF��D�@��S� \�;APKPR� C�G�
D ;EN?CLO�O�S_MCP� d��
�D��E� �3@M�C�^���_MG9A�C�POгq0��BRK�NOL�� ��PR� _LI��1���J �P B������^��Dg��6/%nQ2"8�����!�� ��p�]��'j�#PATH�'�!�#�!u�h�#�@Ұ�CNu0�CAB�@�INFH�UC����0C��UM8Y���C2���E]�3:j�3: �@P�AYLOA�J2=Lk�R_AN(�t3�L��~9z1n9�1�R_F2LSHR&A�4LO41�73�7>3ACRL_�A5��07f4��H��E��$H�&BFLEX�BC�JH�� :U�g���WGnDj�`����s���F1nA �E�G��������� � RE
��.�@�R�d� v������X�T�������@h������mA��T5g�QX�0����CT}X ���e~X	-? C L:^gy��	|"}J�� � �0����l�AT�F�6��ELWP �u��J� �JE�C�TR1�ATNPF��v�HAND_V�B�RBA���$� $I`F2�nX ���SW)�_s���O $$M�0�R��h��x��Pk�"��A@��k0������A����A�A����T���D�D�P� G��T�ST�\��\�N�DY�=� ��ƅ|00�7nA�7�1@m7��+d�@x`�P7% @%I%R%[%d%m%v"`s!� ^�CD�"}�xY�q��ASYM�%�P� �&װ��-�1�/_SH�7 4
-���/�*?<?N?`?r3J�y<* �:J�@��9�D_�VI���q��V_UNI�3���c�1J��Ų�Ų�<ɴ�5 ִ���=���9* OO�Mņc3D;C�$H���1�(�{�ENL��DI�vCO��q|!|��� �`
͂I��A.!�3���@�e���8��pC���Q��o � @�ME?Q�"p��J�g�T��P�T �Lp� ѝ � .��8�,�T.��� $DUMM�Y1�a$PS_6�@RF�@  � s�m��LA� YP9c��� �$GLB_Ta��Ũ�Г�C�&P�q��� X,��!�ST��SBR�� M21_V��8�$SV_ER�0O��p���CL����A�XPO��w�wpO�� �� D ��OB��sLO� I�6��\Ӧ�6���qSYS�6�ADR�qw��T�CH�� � ,xI`/�0W_NA�Ac��\uSR!?�l `��R p��僆�閂�塇�� ���㿉'��'��'� �9�S�.�9�w�ECX� �"��e��������|0�|!XSCRELj:��(�� ST~F)�}��D��{����p_�pA9�� T,	����q� �P�B�q�A��OʐKIS�q���| ;UE��� ��!����S*��qRSM_����UNEXCE1P���{�S_�Ѵ0�3	73uC�OU?P�v 1-�UE�����\PROGM�pF�L�q$CU	�P�Ob� P�I_�H>� � 8(A� _HEB�� ��?RY ?��d�p�Ab�jүOUS�@� � @��'�_$BUTT$Ry�>�!COLUM#�ŞVSERV�s�P�ANE�p9����N� GEU�q_ F� ~��)$HELPe%^��ETER)�' (�(2��(p�)p�)�0��)8��)@�t IN� �� NS �p��1q�@  ��L%LN��� ���w!_e"�$HB0�pTEX�sM0A1���adRELVPDPl�as0E5p3MV3?,�5S3�tq2�шc��USRVIE�W9�� <���U:�@�NFI�p�0�FOCU$��0PR�I[pmc�K��0T�RIP��m�U9N����� ��B���WARN��� S�RTOL���	 t5QV O��ORNVG'RAU:YDTnI����VI����(<��yPATH�2y�CACH9cLOG�G�ALIM���C6Px���5gHOST��!�¥R_OgBOT��QIM�G ��S{РpU �B����H���0VCPU_�AVAIL���AE5X�D!�PMT�G~R�G{�N�``a�@�bՕ9�2�a�Ev��^p$BACKL�AS�@Aq�Ab:���  ��C7eV3@_$TOOL��$�A�_JMP� �<�T �$SS��Yt}�r VSHIFCP���P%�y��� �j RjhsPOSURz�sW��RADI�1�d�_�ӡe��q�P�����dLU��$�OUTPUT_BM�QmPIM����`�`����cTIL�gSCO�b�cC��d1B �f1B�g1Bv1Bw1B"x�D��te~}R�W"�Pbߠ���B���DJUUA8!d��WAITx�B�U�%pNEa��YB�O: �� c$x����SB!�wTPER1NECQ�+�?�'�� O���S1R�Y@g��c<��$�B���M��7!���b\఺@�Q�OP�JM�AS� _DO��
��T}�D@ m���0|}��DELAY���JO� !���ԣ&� �s�0���`��QO�\�Y_�A�\�v��c�A|h$�? r �ZABC��� ��P���C�0
� �$�$C�P;P����ё{вpڐƐVI�RT�1ϟ�ABS�a�1 ��� < ݑ'�9�K�]�o� ��������ɯۯ��� �#�5�G�Y�k�}��� ����ſ׿����� 1�C�U�g�yϋϝϯ� ��������	��-�?� Q�c�u߇ߙ߽߫��� ������)�;�J� �>��AXLMT=PJ���  �\�IqNe�w�[�PRErP�1Pj�����LAR�MRECOV ��婀F }�ݑdJ��!�3�E�S����v���������, �
"���V�NGXA ��	 =#��
+ �PPLIMCX?��Handl�ingTool �l 
V7.7�0P/53 ���
�0_SWq�
F�0�� 154�2��v�7DA�7~ ��
e��{:	lNone��m 2P����T�GX	�Z�P_�!V��Qu�6U�TO��;@k��Q0HGAPON�d��zQ1U
@D 1��� ����S�Q0�`Q 1�� � �������	�6/G%��\#֒�ܒ �`+$�H%�A*HTTHKYU/ג/*/</ N/�/�/�/2?�/? ? >?D?V?h?z?�?�?�? �?�?.O�?
OO:O@O ROdOvO�O�O�O�O�O *_�O__6_<_N_`_ r_�_�_�_�_�_&o�_ oo2o8oJo\ono�o �o�o�o�o"�o�o .4FXj|�� ������*�0� B�T�f�x��������� �����&�,�>�P� b�t������������ ��"�(�:�L�^�p� ���������ܯ� � �$�6�H�Z�l�~��� �����ؿ���� όZ,�TO BTDO_CLEAN�|4��NM  ����*�<�N���_DSPDRYRL���HI`��@�� ����������(�:��L�^�p����MA�X? ��Z������X�ā��6PLU�GG��ǮRPRUCs�B������ĝ��O�|�4SEGFzKX�j�u��� �ϼ�������<�o�LAP�߬�n#Xj |��������0uTOTA�L����uUSENU��� �ȋ����RG_STRI�NG 1r
��MkS2�
�_ITEM1�  n2��/ !/3/E/W/i/{/�/�/ �/�/�/�/�/??/?�A?I/O S�IGNAL��Tryout M�ode�Inp��0Simulat{ed�Out�<OVERR�п = 100�In cycl�5��Prog A�bor�3�}4S�tatus�	H�eartbeat��MH FauylGCAler$I T?BOTOfOxO�O�O�O8�O�O�O ��� ����O5_G_Y_k_}_ �_�_�_�_�_�_�_o�o1oCoUogoyo�OWORx���a%_�o�o �o�o!3EWi {�������8��/�PO�A U��k>�x��������� ҏ�����,�>�P� b�t���������ΟP�DEVX���l�� � 2�D�V�h�z������� ¯ԯ���
��.�@��R�d�v�PALT ]���ow�ſ׿��� ��1�C�U�g�yϋ� �ϯ���������	ߋ�GRI���Aѵ�� i�{ߍߟ߱������� ����/�A�S�e�w� ����/�iR]�� Y߿���1�C�U�g� y����������������	-?Q��PREG��� ��c�� ���/AS ew��������W=�$ARG_��`D ?	����8!� � 	$W6	+[L(]L'�W7m)�+ SBN_CON?FIG 8+�1��2�!CII_SAVE  W4��!�"+ TCEL�LSETUP �8*%  OME�_IOW=W<%M�OV_H� ??R�EP��R?%&UTOoBACK� �-�FRA:\�w Y?w� '�`�0w�?�: n(w�?O2O)O8;OhO�4���nO�O �O�O�O�O�Ow�O_ ._@_R_d_v__�_�_ �_�_�_�_o�_*o<o No`oro�oo�o�o�o��o�o��  ��1_q3_\ATB�CKCTL.TM�P XLED.GIFas��f8WINI��w�%�k3MESSAG� �q�!@ �{ODEC_D� �&�6�xO����k3PAUSU�!��8+ ((O ;"U�g�Q���u����� Ϗ��ߏ��)��M��;�q��0�:�TSK�  @��?�n0UgPDT�p�wd��
�XIS� UNT�E 2
8%�# � 	��'�R!�O� :�s�^���������˯���MET��2��Pܯ5�دY���S�CRDCFG 1�8%B! ��%�"N���Ŀֿ� ��ϛ?�?��T�f�x� �ϜϮ����=���� �,�>�P߻���'#q1�GR��ސ���7pN5A07+	q4�ַ_ED�p1��
� �%-=pED�T-y�/:	�-�����$0-q3��w
�n"dOw����2 V�.;|���r�	�J��8
�y��ED3���g�����C����/�ED4��V�z�����8R����ED5B�������ewED6��S���/8�	ED7�B��f���>/��ECD8./�/2���pw/�/Q/c/ED9�/�/??�/��?�?�/?CR����?�?-��?(O�?�;����NO�_DEL�ߩ�GE?_UNUSE�ߧ��LAL_OUT �@�t��WD_ABOR�p�N���@ITR_RTN�w=��LNONS4��v��q�ECAM_PARAM 1���
 8
SO�NY XC-56� 2345678�90�� ��p �@���?�H�( А>Z=�F�]Uu�f^@UHR5SSp=�vѕ_�_R57�_�UAffjZ@O0o Bo>OfoxoSo�o�o�o �o�o�o�o>P��zCE_RIA_UIޘ�PF|������=��q$SG�P 1@���~u���#��{C�I�D�F�PC�pCe F�(F�SPC8F�e@F�HF���CXF�U`F�hF�pF�x>�_�� C�F�����F�����ɏӆ=�jQ�PHE�0ONFI�G�O�G_PRI 1������}� H�Z�l�~����������KPAUSPO�S 1-[ , E����,��P�:� L���p��������ʯ����:�ВO|�����R�NDET�_V����C2r1KV���r��l���PVc 7ܿ�y
 y�￷q)�;��<�'� ���;Y�k��Ϗϡϳ� �������T��1�C� ��g�yߋ��߯����� ,���	��t�?�Q�c�����y�GRP 2����r i�y�I�O ���Q�w >�F�X�j�|���lF�}�TR����'�
�E�_MOR����| �� 	 	,P> tb���s����񒒺A?�큠��pK(��R��PV���j�a�-�/ A�tp����u�ȵtb�wi��hvPD�BX� \���
mc�:cpmidbg�HO#:��q����p�U/ #  ��p�F�����/d*ܷp+w/C/�/&e)�88~(g�/+?�-E~(f?s?)�u?~�DEF ���C)�b0buf.txt�?-�?� �_MC��!�� �d(,EC��"���VW�{�Cz  B�q B���FB�8�B���~C� Cޢ�D3�u�z�q Dzl'D:��"DrBENN�EA7EV��ߓMF�pgF=�C�F�e,G����Gp��G��/��yjT	F�$���4m��p(T~*�p�p�G0�VT3P9���A/  TRy�{D�VPa  EY��E� F*� �F|�G$ˀF[ߺ GR�k^Gl���G��G���&H��G֟��H���C���  >�33 s��A�  n�q�@�B5Y�Udu��A��t=L��<#�
4�1�o'��BRSMOFST� �>�rIT1><@DE %�l"� 
 a�q;�` � 0o*oNTES�T�2#_oksR�r&(\�#^FCPA�[�B��aoBՁy�B�@�x���SN1uT�_�0PROG Ċfr%�?��vIN�USER�铄vK�EY_TBL  �7��Z@ �	
��� !"�#$%&'()*�+,-./��:;�<=>?@ABC��0GHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾���������͓��������������������������������������������������?������ё�p�LCK�|��s�pS�TAT�s_AU�TO_DO  ���F�INDT_ENB;�w�R�aY�K�sT2���uSTO���~�R�TRL�pLE�TE�� ޚ_S�CREEN �FJkcsc �	R�UϐMMEN�U 1'FI  <�|�l��K� u����㇯��毽�ϯ ���R�)�;�a��� q���п�����ݿ� �N�%�7τ�[�mϺ� �ϣ��������8�� !�n�E�W�}߶ߍߟ� ������"����1�j� A�S��w������ ������T�+�=��� a�s����������� ��>'M�]o ������:�#pG+�_MA�NUALӟ��DB;COu�RIG��$��DBNUMLIMҸ�,Au
�PXWORK 1(FK�o/-/<oN/`/r+�TB_� )�}��Y@$�_AW+AY��AG�Pr9=�`�&_AL�=���"�YҐ��p�_�0 1*�k , 

.:/�d2?o?��6� Mt�IZ`�,@|`�3ONTIM��t��6�)
��u3MOTNEN�D�4RECOR/D 10FKUB)O�1�O�?A-O�k�" kO}O�O�O8H�O�O?O �OcO_*_<_�O�Or_ �O�__�_�_�_�_�_ o�_8o�_\ono�o�o o�o%o�oIo�o" 4�oX�o|�o�� ��E�i��B� T�f�x�������/� �������>�)�7� t��0p.u�����-�� ۟͟�����N�`�ϟ ��o����)�;��� ���8���\�˯ݯ�� ��;�Q�ڿI���m���4�F�X��"TOL�ERENC�$B��	2� L�ͰCS_CFG 1 ;�x7dMC:\���L%04d.C�SVY�0c��x3A� ��CH�z0�_?x>�Gߠ}<��R�C_OUT 2�+-0z?��SGN� 3�%�2��#��12-AU�G-25 17:�24�O27�-MAY��4:3�8�]� Z��t�����x>�з�p�a�m��PJ�P��k�VERS�ION ���V2.0.11�~;EFLOGIC� 14�+ 	�TP��P��p�PROG_ENB�/\B��ULS�7 �&�p�_WRSTJ�N�0��2�$EMO�_OPT_SL �?	�%]�
 	�R575x3?�7�4D�6E�7E�50i�d�o�2E�T��j�>"�TO  .��l��k�V_�0EX��d�5 PATHw A��A\���M_~;ICT�!F�� 5 7�$`��eg��}ST?BF_TTS�8���E�3`���M�AU���2MSW��6 9��}<tТ�7�*!��]lR��v�����DSBL_FAULy��8�/�3!GPMS�K��2TDIAG� 9���`����1234567890x'S�lP���/�/�/�/?? %?7?I?[?m??�?�?��?�?�?L#@PV/ ��"�/��  2OXOjO|O�O�O�O�O �O�O�O__0_B_T_8f_8Lx�UMP$�I�3 .�QTR>;#��_�PPME��_Y�_TEMP��ÈÓ3��4���TUN�I	�w�YN_BR�K :��x�EMGDI_STA	����GeNC2_SC/R ;7k�/�o �o�o�o�6�o�o 02r�ncUa1<yo+O�|����lbTt=7k�Q����� �o>�P�b�t������� ��Ώ�����(�:� L�^�p������� Oǟ ٟ�0�,���+�=� O�a�s���������ͯ ߯���'�9�K�]� o���������ɿ�� ���#�5�G�Y�k�}� �ϡϳ���������� �1�C�U�g�yߋߝ� ׿��������	��-� ?�Q�c�u����� ��������)�;�M� _�q����ߧ������� ��%7I[m ������� !3EW��{� ������// //A/S/e/w/�/�/�/ �/�/�/�/??+?=? wa?s?�?�?�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O�O�O �O_K?5_G_Y_k_}_ �_�_�_�_�_�_�_o o1oCoUogoyo�o�o��o�wETMODE� 1>'Ufq� ���oGwR�ROR_PROG7 %�j%���H�wTABLE  �k1_����j�RRSEV_NU�M �b  ���a�pq_AU�TO_ENB  q��cZt_NO�q� ?�k�a�r�  *�6��6��6��6��p+5�O�a�s��HIS�sXq�`��_ALM 1@.�k ���6�6p+t�����&�8��J�x�_�r�  ��k4��b���`TC�P_VER !��j!6Z�$EXTLOG_REQ��s���SIZ�~ܔTOL  Xq�Dz���=#�=
ޒ_BWDo�%���vQ���_DI?� A'U��dXq< r[�STEPg�y�|�`��OP_DO���$�pFDR_C�FG B����?ZpA   >π  @��أEATURE C'U�Q��aHa�ndlingTo�ol 7� 5\r�bEngli�sh Dicti�onary=�60�5.AA V�isS� Mast�er0�>�0iB/�a�nalog I�/O7�>�PRIN�a�uto Sof�tware Up�date  B/�16��matic Backup;��duct��g�round Ed�its�  D p�rCamer�a��F��1
P��ell��ʱ7i�n�ommj�sh��8�8\hi%�cyo��=�ct\h%�ޡ�pane6� R� J8%�tyle select>�7\im�on߱j��onitor<�h�73x�ntr5�R�eliab��<�0�y�Diagn#os����:�
�����ual Chec�k Safety_ UIF z�1E��hanced Rob Serv���q oͰ�UseOr Fr�>�A��E�xt. DIOm ��fi�� #��=�end�Err���L��\�6`�[�r䀰C� @�:�IF �OFCTN /Menu��v��>��g H��FTP ;Inp�fac��?��6\aGذp�l�k Exc	�g�5�Y�High-S�pe�SkiƳ � ��!)���G�mm�unic��ons�>� M-��Houqr��p���R Hx������conn��2z=�(�Incr���strΰi�<�
�TEKARE�L Cmd. L���ua��pV�s�R�un-Ti4�EnvU� "Tq�z�m�u+��s��S/Wɲ�
 �Licen�se��'� L��o�gBook(Sy�o�m)��oad�MACROs,~��/Offse��/art ��HG�R�\ap`�Mec�hStop Pr�ot��d� \h6�4��ie�Shif8��9��MixЂ�ܾ���CVL��od�e Switchn��c.p �Mo�����.� 72l_d����g'�l�!��?ulti-T��⳺��!W�Pos��RGegio���d#�}Pr�t Funb���II)��Nu�mЊ�d� .co�m12� Adju��:�41\LZ� �J85P�ktat�u<�mm7$�R�DM�otN�scwoveW� 44W������uestO 7nu`��oG�܍�<�.fd��SN�PX b�⊸50yS�[�LibrV�N'"Lo,� S��Pa찠�Et�s in VCC%Ma0�ѣ� ����Z£�/I����T�MILIB��7:eP��Accٰᵞ�TPTX"��0;iCeeln��Ar�e4��8�O9��Unexce{pt�motn��  U�) -�7�N𴰌f�� 
��a& �t�Ha&SP CSXC9�����%[�3�{ pI We�4'�^ \�$vr��	ҷmenS  N�i�P^�a �
7Gr�id�play �����6pŴ��0,&�LRl���2���%�K�Ascii��l���7�ӗ�st1P�at����OR�yqc���� ori���� M���ata�qug�c���[�,�0�-���RLEam���$5��HMI �De�(��� 7����C�߇�	 ��a�ssword?�LD% � p����7�"A �YELLOW� BO�4Arc�V vis����IF�5t��OpA�;�s�^��sp 2۰a���po� ����Ta1���2� �HT�І@�xy�"V'���l�lig� !Q@@�� �!0JPN �ARCPSU P�R\<�9��O�L?@Sup�Bfi	l�0Z�2C!uQ^�l�cro�mS�L4o EST�SS?@]ee�tex^� J ��Qo��t��ssaIg��@�mP�P���]�!	62_�Vir�t���9�z�1st�dpn6���SHA�D�@MOVE T�F�MOS O��4�5get_v�ar fails! ��o`%�AE۰��� Hold Bu�s$$CVIS U�PDATE IRTORCHMA@$��iWELDT�S� st�Q�a: R�741-�ou�`b���62�!BACK�GROUND E�DIT Sb 26�.f� EPTCD� CAN CRA�SH FRVR �A/R@�cCra�.�s 2-D��r���$FNO NO�T R�POREDU �p .pJUPO>0� QUICK�`O�P FLEN�L�oc���bTIMQ�V8�FPLN: �wW��plT�FMD� DEVICE �ASSERT W?IT 823`�s��ANTqACCES�S M��JoQ�ui��<�|r��x�U�SBU-�t & �remov��,S?MB NUL	@lq?ER FIXG��HIN]aOL�pM�O OPT 23�g `OST?@wD�U h�p�dAddf�ad.е@io �� AMpP�pWOR�D.$apO�IN�;�50�aP:fi�x CPMO-0�46 issue� 16��J`qO-�P130��TE�S�dSET VARIABLES^`x����c3D m��view d(ML�W�ea��8 b.�?of FD ������Px OS-1�44 ��h s �c
p�t�s ��lo �� �h�WAp��3 CN�T0 T iLB��T�Im��Z�ca� mq� POT:W�hen��ews�STY M120a��t��pt|ado /GET_�� �,�VMGR qAWpA�@C�a Pq@�C@��ͱ�� C�@� EL�ECT?�L<�IN?G IMPRPQx��RY�\`s�PROG�RAMOP�@� IP�E:STARTU^�AIN-l�  =ga�SCII�`���OF LO��PT�TB: N �ML�K4me0��:��moW�all�pR�L�]8l`Tor��AH�`��yS1QP�th�p}n�P ch -рp� yTU@Rtou��>5�iRCal��Sign� P��xU�Thresh12�3$W�Hj� : �MSG_P4�\@e�r  ap�G�A�zero5 ���@/ 6tc�d:��U@���2D� rc�O3ME�p�ON�`f�| 0;ASREG:wV�^�őHt˳KANJ�Iصno̐0Аc�@��n d�1�QTE�Q�INISITA?LIZATIpD�Acwe��� =�dr\���D�c��minim9 rec0ˡ�c@����mU�ro  i!C�dϰ=�i��(�{���vdw�� 0iqB�Ѓ���w u-Ѷmse$SY�`M�-��q�#%�bW�l�u��d�Re�eÂ1|T���m t06�0�Warnő@�בB�ox fo�Pse~qPVERWRI�`҈�S�¿�F��up~�de-relc0�d"�������őbe�twe��IND �*��igE sn�ap��usősp܇�FTPDT�DO��TqHANDL �  ��d���D4�n�  D=�����operabil��0  H5�[�:� H5�0l��ܲ5�1�!����mp�qs_  J52��O�p�FA�P_�^aV7.� )U��`GTH�pEi�sݐ�0��mq����ne-Rema�rkE�� RM-� tpqtQfPA�TH SA\`LO�OS��[F�0fig� - GLA e#li�з���p'�ڤ|d �!Ether���� Trac�� H55�W@r}7O� 2
PE�H��>�80n�P l\0RQ:��Ɛd|�y���it �P�p��Pa�y�1[2]��
�X^e1: g*�s���dowDt[ �@I�S ���EMCHK EXCE|�1H�OMF +���qh��PnHPZ�P�qB ��Ĵ��Xr�8�0 �r��c?��e A���E�Fal1�ala�rm�� V��IRx`[��v�1�r��a3opX� ck��6pr � "y��@x������Stud>�̚`b fp��: U�0BUG?��2��DUpPET<���� ��S�EXPANS�I��DIG+�KPO� ��dCCRG �EN��CEMEN�T �pHM��K ����pH GUNC�HG�`�EXTEPpP�cғaS� 0q������ORYLE�AK?��4��pLC WRDN R1�qO'�
��SPEn����G[�V *�|!MpU�=�7�SGRIH�A�@�0\t��M�C ETH� ��S�Uh��p 8Y��PENS�`N�P8�[`<0a��BROW�pR��RMV ADD ���rA�DC��pT�3 ALAcP 2���-�VGN EARLY�b&�����8wr�!LAY{�8�O SPD��[PHM#�S "T1�0TOGUCHi��Ї�F���JaY�y�5 _ERR�ORF DE SA�/<@WRO5�CU�RS� i�I�N �np| @�[!-158x�G���RSR �`BTqU��7@�6T�"F7�"�s�%1�%�u�@!B� SY RU�NN4���9�p@�BoRKCTARO�bdP �@�`AX�`���PƐ��@��IS�SU/3�C$pTS�I�1KWCIPSAFETY C(7ECK|�59=#qA 4�w0���=�� \!7TWD�R41ǱC!�INV-�D ZO�P��R24;%z21DUAL6��ӁC!S�FT�E� b���!0?NDEX F� �%� X��%UF�BP���h21!�4RVO_117 A	pTg�q �PT�@�FAL"�TP247�Rt\rSQP[A�HIG� �CC��SNPXF MM�!4�@��t���V>�\��2`�DETEC `p@�� "RUK2�PuOS5��Y�6L��G�� ��vWT� �� �9691U� ROP�P�P BFITP43MS�qgkϑ@�RCOPYG6IAL_�[ T�@4K�`�6IA"GC�U� i�� �`A SIZEO 674�`O�7��-\0�!F_RO���D�CP PA��pAgNUC؀S�IL�'.pc` �`RE�s���ple��  g�tpa� �`
��a����\r�b���utl�a}p�`sn	p'�1{p vKt�21up|Kpcirf�b� JqslDq�htpx1!spnqgi��Cxkey�}�)qgvpm0zp�|u�su!ug-�.vr*����b��s�]��0��$q���!! j9�21p��pl.C�oll	�Skip��y�R��J��*�3�d� ��i�q�� (��, x� �Ar v���.�]~���>w2�1\at*`7 "�KF�Q�,����\twptc��"TCX��m1�}e�pkmai�n�;�setskck0|ate�m�s�Fș�郣�7���KAڱ�U2 Sp��FCCTN���0ЀpJ���ڌgՀ7��AREAL�������7A�@����)�f�)q*`8I��8O����h�D�9�I�9Q�pz�k���r>p"KRCF��s��ڢctme "�CTMEO�Z�أrcf��p|�(�!����g�pcfcstm8T���,�cdt���� +�s��rpb��ٖp󖦅73�P��p=�� ��� J�$��q(K<�� N�p�� m�p'�]�p����?� b÷�pr�c���U�� �rp���9���,��� Y� ��qv�_���p��� ���̲�q[�й���V��52Zd�C� �uh Set
 � ��� ���J	p	  � r\tq_zm�oveo׹�fin{de�ornt�`��Ѽ{4�p�L�p\ofndrٙ! 4���r�tcpmate��T��M����0�R638 R51Q7˂)���(��aDqP�	�t(q��m�%�����B�99��8�pp�0,�i���p�PM��)��etguid "�GUI@�y�V���s�pe�)q.�tm_mqo������refB����a��)�)q��lo�g�P��prmpA����va�(V� �����������	��/mask��Gq���sk Excha�nge����2H5[41%93*0%Fc�96%0&9%"B5)p?2��1��uN��v�m�x�� ��0I�0k��t� "�1£�}���H����Y�dsukch�P�sDi��yIm"�v҂8|@�&�887 (G!>]�isplaT%� �RƠ]�9%�x9 p��"*`2I�2O��+t
9 c�D�@x�� ar� 9&�߳(1sca82��*m�scrL�BsX8trld��S=���9(��p8A$ayl|.��`nfirm2#b'78ڊ��A�  K���@!��{8B�3�I�3�/]Ei�plcf "PL�?�D�pfca0�8\`�A����D�Bov�?�Yinim�~V.avp"&aA�r6�A���Shape G�enerat��IIDQ��74ڈ�r�R (�]p�(�p�a��^|����K��enuu�\�hD`n�HMN8:A�;cil\D`<`�sug?cia�nue �Bshfi���fhi` �Ofd�!��tm�?���fh�a1vY�$|2��o�k�a3<�io#dsm;jenR��>7mensub~~}�`fh� �w�$yseQ��w2�rc�MSfhst0H�kc�Q�6d��lbdetbo�k�gk%E^fg8��
p���	akadspweb��Vo�x�����S���G�:b201��Y|�3�����!4��9d�5��"'e|�il��@�����[,��HA���� (CalP�,q�_a�ca=�_	W@�4�6�;�6�ϛ�ţU�mt��LMT�ͽ�et@��ALj�-�몶��7ţmc��K8ån�sv�3���� Q����c_�@i�~Y��joi@�ٟ��F Y<��_trc@:]�o����c�������0�@���4�}UCenter F5��1_�20\0{��ɚ&@)¨*4�/p�5�7;��7�q/�� "F ���.����;%�4�@�����ٹ�.��qp����W�a��g �  uxra�p?axrmrf�oG��x��"&K�/'tur_bsped�T��\��W015�P2�����s)��(��ya�_��F�⦯K8��P�k9�7Т�|�$�1.�8�K�78���'�ts�p���1?"���gglfmԏy�st��&�R�O�*�vAr����� vQ����@a���Y�| p�shim��P�Pi�m (xTool)T�6������ ���Ale��]q�`�	�5 B�fx@a? "TPSH�s�'pe��FLEX ���'1�5 b�R�R�r�%� l�rE^P5 2Aѐp�����padqG�DQ��5 ]�8K{ �A4@DQ�_��7!	��1�s7�!/�95��+�1q�vl "DQVL�	d�$dq�I�I�&�c3c  �H552_�-121� !dAAViMS-20QpaE0�TUP s��J545o�i061�6?0� VCA�M @RCLI=O�#R6m0� ;dq�0MSC{c�2�P�#STYLk r9 vu128@�+��0NRE/#�0S�CHSDCS�U rmal�0O�RSR c�u10�4��EIOC� 3�Q�0542 ���@SET Ea[sy�0J5y0Uk`�(i07y0��MOASK ��27#�>�0HOCO )�5B�3�Ci22W�fik.5B0 8֠#u1U0�p5539_F�A"N�ORMLCH�KK5OPLGQf�ii103�0�M@H�CR�M@C�0aAf��B6��i154wEMDSW�BuQi@����137��B0�Av`�@7@P+��C7 ��r5B53�5B7  <A��B5�SPRS�T 77a�F�RDM  J98�9�0�1��-0930��R�PSNBA u�hQ�0HLBGESM<�PTDSPVC#si1q2V0-0TCP��?TMIL��P�PAC k987��QPTX{��PEL�N�c�B97�UoECK L�88-`�FRM ��� �1OR 8�0I�PL+UCSXC �e\sw�0CVVYF�QTP�Ad�@���6Orob�0G�y`�I�Г5I�PGSns-08�%`���P��7eR6�63�pse0Q523 "rkey%R�1K5R696{g5k1 �a.A53�U֛01 ~`sh31 �a��4A6%`�AA7G5 t� �0�`6ca=l�`CTOP[�A��0>pc80 sl{er�@PRXY�5�7p0v885 r�ec;QOL�0L4S�}� qe�0LCM� h��lPETSS���%R6��`�PCPsE ��PVRC��t�bNL�eU00'2 u�3�p6� <p�r7 �at�q�@$�R�1�e�4�m��5 > W\0U02^"@se CI�3sU�K�4 822rK�5� p��q�P(Wai(��`R�o<�3v@��\y�VU046Po
&��3 �"��435��C6 .��q10�A1قy4�Eۀ5 ac��~ق7 "MCR`�S61oe�4�AmH��65 96J�	�6���PT�68Ǉ�qpMa�73SuG�770�qipM�̂83�5k�4�"<��pw��pk��8�Uk�9����q9�0 w�s��1�9�"@��95 f�u9�7�5U15P����1c01w��vFU1M����H�1qP���7 ����8OP b�PU)1�@=!BA�1OR$�	1AQw�6�P��?5 16 (L��`�o"�NP�푡Pt\bu<�1�`�z���s���`��!@bbf`��m0dǠ�fU1U0Obox\�`�1��68,�1P��58���59`69��60ק����p'��6 BBOX �6�7�u'���pschme�71[�72g�?6 setu�����\��p����offs�H�93K5ð�b?�2)�btas�@۰���21�219�Pl%d��2�`��2q��:��2!@xcdg1��8o5�9 ���2&U0li�E�23�Ep"@�55P ��� =�<��5�p�4k�3 or�^Rk��pro'qk�63 y��i�7 �i9[�R$��A����2� P Eoq��6 �very,��9 ��i��ʃ5q� ���8��5�P ��`���5��971"��3���5��e��!@ecj�aO�
@��i��`���	pK�q�ƀp�p�80������6 ��ҿ7 629 @@U�5�panagH�5,����57��5��*`h�a��7>�57���Մ582 4�5�y�ĕ5��o�i���"�XRM@?�2 C�  �=�3 	��K	=�4��99#�6�@�y��@�y�u@d�6AP\ac�ׂ6��e�y��0ĕ6ҡPvt���6��"A+CS��7{�6E�_�0�qc�0�q�\�9��sv�`ANRS[ e�r� vs!��h���Norch�ma��� � =�M�a!�!�� 39 �J59!�598 _J681 !�7e�`J6Q�W%!��c�!�L�te,t�s&!�`�P�#��A��� �$�IF!�AARCRNt�1 H��a�o349�:�\9�cp���P���s8�FA!�H�597��92!�L�SE�#]�[!���t�mk]�4`60�A�	 ��F��t�1%�0!�&!��or!�S961!� �!�k Z�x/0i�!�9��?���f_ �!]� !�� !��4��)0i���(��tm��]�>�R�h����A� "TMA`�&��y��in_!��A����Mp�!��&����etd�2���&!�����moveto���%��?�9�mmonitrD��&!�x� �Tonst,"��a D"YDP���^Q�! para�HI���ame]�C?ontrol8�W�,@!�43`�0@^��25 R0�588�P0�`��t�]��� (PP�eter�"!�,������R,$ �"L�QmB�;33�� `\ �E/93�ap����e�2� m2�ol_adj.f]�T=p� F�2Adjus�tA� `��1�8BZ1&A�J (�2��e �3�$2 ��e02j�2\P�E5�`*C,�adFA�DA�
�� .@t� �4��m10s>OPGj@��O+B��p�	!	��1�#8�`��^PI��!�ae�1aBi�3���N5�3 H]�(D�r,�ol 4Y,4 Q%r��ᩢbLaq�r� �5� !�.<r �E}C!������vC3S�d`!�fi��PFI�`NyXsltpalx�_�Ztpts�TSRN�[�{S,�pf`
 sw��\� ��J	�!�	   ��J�-RServo Gor������򑠂u'j��bT��fD[��އ�j670g "SVG/`Q�eQ%��aA2py "CO00qX�, 0��o�f�sgn "FSG� Q"7P.�`s9f��XaPSW�
fB��A�e	!sgatu�6p!�e��asgt=p!TPDR0o�j�bs�19�79o3��(sP��t,��`GATbOsp!�[sr*>�bsgk95*��W�Yq?�ftdL�ߐ�������rtdf�l\!�Jځsmc�hh/b�tdmen8�2I%�mkpd�1����xhk�wmvb�󈄐ku2�f��mklw�0���fsclini/)u,�Oldvr�"�v�1 �X�9�J�,Q����`�aaut�p�7A�S�8��1re�sub�'P!�Nt9�aZq����b4Au��Muh�ĥ�hk_kvP�Y  >�Yq1��P�H1�ف�tol.p1�i 1�7�H �1�G��`1��sev ��1�g�u 1�w�K 1�x���`1�kksk� Y1���, 1����1�.Ƿtch1�q*�$� 1��p1���E ���uk݀��$�v�1�'�Yp�1�7�H 1�G��cl�.�d�!�t�1�F�\	j1�J�r�a���1��v�VL!�Ĺ1�gtsgvaٴ1��q����1�Ƹsg1�ex��Y1��0����p9r1�7�cre1��3
I1�&�571�6�du1��bf4p�A�π����B��E�%��a.Af1��B���� �c�Sche��T���Ho�44� 8P1��%���S!��d+�1� 2  �H� 1��	�Ktb\q��tp��0b0l� ��1��D�+�trackin ��0����P����enc�01�����q�i�K!1�������altst� ��E�б�vr��1�e��P���ם0���41�sb�a�CVers1�ll�Bk��!S� �(Qv�"(V��Bel=U1I��,6}�baaUH0�1�u��ssT`E `�
d����b0k�j05��sb��9 I� ����9�F� ���B���en���C��(QD?evices��:��K������41�86 c(O�P�q�es 6)�P��aU$zA�o�\p3k!��j1�p
b��@�Zaopn������|�1�#pc������o`��glfm_���V�`��&���V�sc���a���цvropio�@q��E$1��A�,�1�)@�����8�18�CNEM��m�p��J� ���! (;NE�ump��z��� 1�F��1nm�n�6��SeD1�42m<��T`MPTP�RA�� 61emocol���33mpΐ���<�"�j536�A1�7uch$�ns�0p1���J5p���$S�32T�41�ngP�% !6p1%	P�3y6�d1THTK�1�Dq��0\etth��THS�sJ11*�0�1�hpgio "PGIO"PEp�vCthwkf?F�Mc��MHC5�4�8�52�V1�xAmLP��q57c�� �F�51/�F
Ttsn��SNSx�����A�1�8V�Aq?SA[QuiAf��Q��*�xAp@ѐt/uD�A�M0�6X5  Ѥ��B^P�ٙ(�2� 	��Ѹ�dQ!�`��1R�J؀E�N�y�1� �s�J��1�ipc��x�ݥ` "ctsk�e1*�`�R2k' ��!�p�a��!�acc�0op�4pC
p���R630��aX�)pp��tt�!Q) "q�u\ �:DJ3��r���paachZ@ACCH��dOfw`�4>0�K94D3AO �u3k94���p���q����chflo1 �ST-�v�/Suq��h��fp�A9�st@������w�l��)�sA�chcal2L�^�6�s��@�F�0_�%I�[�vr	r�j|v1�! pai�a�Q�RA��Watecrb@�����56��)L@���5=0(t���}�rnet�!QTy�$ j�5B��xv��ؒj�a�ICSk3o`�\p4�p�t�s���&�1�`�p�w1*��k�ta�`��k�cc����D���cgen^����!cf��C�Ԧsp�E�Кpaw����ؒi�c���O"D���ѱ���q�Fg�!�w��A氂ow��!�R50`�@�3����ư (0�F���/*���5C�q4� �$q��r�x!�]`P��Mp1�Z�55d�A)���ѥ�*/|�aEf؀b����U�a�0i���(���af��|�ep�0��ca߯�����Qh���u���2! ���Line/R�ail T�䷽69ɿ�� (����� FWq�i�0g5OGJ��p8�r8E7��\�9�r�0E	�%��q�53R3=� ���f�aldebu����Rkr���q3�R3RA� ��pg{db DBG2X�@��!
��ۀ�� ��2�2Qҙ% k�Ѹ�ؗ��`��MH_bpe�r Option�c�78���	P� ���`�����Z'h�g�`9�m��ht�_3F�q�mЂ3@k�At��qd8iᏣa9���&�etw��1 Fb��plu� -�._Handl��O�qh��&V!�G�P90�P�7�A�9�Q(Ma ��A����0Uy�0ܟ.�f`138��F�
!� �hH�qE?���x u!? ��O� G�"fhnd? "FHND�!T�&g��wמ#�Ic���lio�#Ce0�/�O�+CLIO�A1��񑑜 45�A9h�C�14�R S�[UR�AR�!J�JO�ELSE��1���";(CAI/OG�Bp%H�$�O \c��G1��Q�55h��e0tcm�ACMI�pa4�d6t�a�0L0�1�1��a�2iomGenu?�qAf3l7pc 1��8��� F�x�e2�dte1+��9dt��|�7eFFd���b�W`Int 1l P�ump Cont$� ����a`1���4 (�A_"�Hl,$����E�!�ha�quy����apa�y���5 �q�r�q�?:Sa�``1PCD��n���e�`Gcndj��Rq�p��a[O�Qѣ�P�Q_����Pa$��� ��2k0�� ��a�Srt���?��Q�Qd�b!o \ � �����	  ���#��� �&���$�J517 (Progra�just�����`�� j$rG0�0���Ds1�j "P�ADJ���FrprOgadjoAup�ppE�A/�v���3�v�`�f�Dp1���j53�9`�- KARE�L Run- �E3nv���! J��#��13���`R0�J#97�!�"6�!�c�!�a�e�2�"������F�(2+�ime (6U1qe�����.jp1klut>��"UTIL@#��\etqm_"MCGR/ڄ H 1����11Cp(�kcmn����Q��J�\��s`ߖ�qq����ex�<M&�q�tr$�f��������tp�pst�s����a Sta�tus�+P�ѩ"H51 e�"v����g�Җ�зPR70( �17�p��W���&��a!戀;%�Q!sHs2���y%�  �STD RSC~�LANGc�5�أ5�prscr�n5��5�֣Y�.v�5�i�5�+�5�ds�blfl5� Diwsab5�lts�5���C5��#5��ӡ��25���le5���aar5�V5��ds5�`�5�U3�l133�`��5��5���t\��"DFLT5��=�w@sbf5�����
M�du�.a�i򹵝��j550.��q P5�5�J��_Ÿ�~5�0 (Adj��nq5�	S5��Y���`5�zq���5�34��ݵM�E�d�q��Vs���Jb!�*�sh5�AP0�5�J#��\a���R a���+պSY�W�M��q�� �C���4�'�p�Sti�PĹR5�7�H|��5�(&���sk��,��RRBT�"�OPTN ��� ���b��K923"��d���03ol��gP1 ���������rcm\pv��57��DPN����K�ccf[�J� I� �K�,�K���J�h�J�o,�I��QI��I�	l��I�s�I��Ӟ����I�ncy.0�UGPDTG�����o�� ��� 3���I"�������iov 2byn����l������Q����
����acc������2��p� 2 ��ɒ��L�R����R������.�a���� ����Q�!�+ -�����������2����������� �v����ex8����	cchW�F24	m�aq! �H㘦w!uTo��s@q�!�汮��Ry&P �n��u-1�82��iag�&Rq �!����5��q
�p��92DP��) �� 6SE>���pi��t�G��
�pg8`%p?�4mon�?z?�?�vr���?Dgse /��f�aE4! 7�e�A ������y�F3�b�%�R823�%lA�c ��E4	R.���5��Oslk9�Ur���*FP26E48ÚsT&edg%�O� �GVTDG"%*s1l3F�_sl��_�Z|`s�_�[�1�_�[filO�\<I�-�6 �X8e��4�U&zK�J5ٲF3m�%5 � �E4	�K�	�O/@���?��tstn�ƕ)pD��)pite ptoo�)pƖMq��p)pEru�lsu)p�v)p^ttl)pjt2.)p�v)p��uiMqtupdc3yc��|vr�P���x�1�����N1���qteq��)p�Ir)p�e��3���o��"�7�@q�4����?cy�r\�dqil5œ)ph��r��l6Ŕ)p�eq��pqA7ŕ)p����Dsw$�,>yxf<�ǖ�]u�Frlk2dq�*��conC ��wcn�vu���bag�tch��pal�ctr���slp|ğ�init0"�4�mnph�z��q����)fя�bT�iu��Ccy�R���Dsv<�H�𿯭�b��s<��d���h%�ߍis��axis0�z�b��=A��Crmled�\��w�ps<Cz���u'304Կ�5���'502�.�3@���� �s��TC��olu�tlF!aam ]T�Box{�I�nw�598�90�`�73CAӦ��� �(�`)� Q!��m�r<�"0� ES�"��sw��`�Y��#F�����@0}�2�\Rc��Yxl� ����q"TL�BX�������olcbx��tԩ�\t�����;� L�x��-!|��- Com�0~��or Cha����Т�Fh!e�OCM R614���B����g ��(��on������nge, P����BT��}v��*��B	�qr<�{xF�p�ak96�� 6�1R_PZ���cr75b0�7� V�h�22h��22~��Ѓ� ��J	�	 �  all<�mreg!"J��?r�W�'�m<�����I�(q��R�m�����>s��5��=A}aF��'�.f ��p¬qaA,�l�qR O Tur����Eu�93 J989h�9 �m�d�"�`� '�Q ���+�i�4�E��N�|��p��P��X���Er��"MLED�B1� ����mk9530ѝ�8՝�����YCSSJ�\�dd�qS���re*��i1p������igr�tM��������">ydk� /*s�$/�*S�<�H�� � �D� |9	��!�!1 C! �  E��  ��# �	�!�"@�؞�H�"  ?����E 8��� �P�<�*�ge�lpq�y�"���'9�9 CP ����$FEAT_IN�DEX  �# ���  � 50ILECO�MP D��=�b1P0�#�U3SETUP2 �Eb5l2��  N �1U3_A�P2BCK 1F~b9  �)�"�?�?  %�?�?� e0�?)Oo5�?UO�? yOO�O�O>O�ObO�O 	_�O-_�OQ_c_�O�_ _�_�_L_�_p_o�_ o;o�__o�_�o�o$o �oHo�o�o~o�o7 I�om�o� �� V�z�!��E�� i�{�
���.�ÏՏd� �������*�S��w� �����<�џ`���� ��+���O�a�🅯� ��8���߯n����'� 9�ȯ]�쯁���"��� F�ۿ�|�Ϡ�5�Ŀ B�k�����ϳ���T� ��x��߮�C���g� y�ߝ�,���P�����tq9�0P�? 2�0*.VR��H��*K�q��w����2�PC�����F'R6:���������T@0@�R���=�|��C0�����*.F�5�����	���� x��$��STM D�MX���E����iPendant? Panel���Hz�j��-��GIF7alMp
���JPG���l���5/��
�ARGNAME.SDT?/��o \S/�/���$�/@/	P�ANEL1�/�/%�o �/?���/2 ?r?7`??/?�?�*3�?�?7�?�?�?HO�*4OzO7hO%O7O��OK%TPEINS�.XML�Oo/:\��O�O�ACusto�m Toolba�r(_��PASS�WORD�O��F�RS:\k_*_ %�Passwor�d Config �_���_�_�_+o��Oo �_so�oo�o8o�o�o no�o'�o�o]�o �z�F�j� ��5��Y�k���� ���B�T��x���� �C�ҏg�������,� ��P���������?� Ο��u����(���ϯ ^�󯂯�)���M�ܯ q������6�˿Z�l� ϐ�%ϴ��[��� ϣϵ�D���h���� ��3���W����ύ�� ��@ߪ���v���/� A���e��߉��*�� N���r�����=��� 6�s����&�����\� ����'��K��o ���4�X�� �#�GY�} ��B�f��� 1/�U/�N/�//�/ >/�/�/t/	?�/-??? �/c?�/�??(?�?L? �?p?�?O�?;O�?_O qO O�O$O�O�OZO�O ~O_�O�OI_�Om_�O f_�_2_�_V_�_�_�_ !o�_EoWo�_{o
o�o .o@o�odo�o�o�o/ �oS�ow��<����p�$FIL�E_DGBCK �1F���p��� ( ��)
SUMMA�RY.DG��|�MD:�[��p�Diag Sum�mary\�iz
C?ONSLOGQ�4��F���ߏn�Con�sole log���h{G�MEMCHECKՏ��J�c���Memory� Datad�lw�� {)O�HAD�OWY�>�P��t��Shadow C?hanges��s�-��)	FTAPҏ?�ΟC�n����mment TB�Dl�lw@=4)�ETHERNET�a��~"����n�E�thernet ���figurat�ion�spV�DCSVRF`�F�X�q��t�%6� ve�rify all�t��s1p�1�DIFFi�O�a���u��%��diff����"�6�1�Կ濎{� ���ϭ�=	9�CHGDE�W�i���u��&ߵ�9��2�����σ� �Ϫߵ�GDM�_�q���u��.�9�FY�3�����ߋ� �߲��GDU�g�y���u��6���UPDATES.U��;��{FRS:\�S���o�Upda�tes List�����PSRBWLOD.CM���|�������PS_ROBOWEL��g\ n�����W� {�	F�j� {�/�S��� /�B/T/�x//�/ +/�/�/a/�/�/?,? �/P?�/t?�??�?9? �?�?o?O�?(O�?!O ^O�?�OO�O�OGO�O kO __�O6_�OZ_l_ �O�__�_C_�_�_y_ o�_oDo�_ho�_�o �o-o�oQo�o�o�o �o@�o9v�) ��_���*�� N��r������7�̏ [�ŏ���&���7�\� 돀������E�ڟi� �����4�ßX��Q� �����A�ï�w�� ��0�B�ѯf������� +���O��s�ݿϩ��>�ͿO�t�Ϙϧ���$FILE_�P�R������������M�DONLY 1F��Ņ� 
 � 5��Y�0�}�=�f�/� ��߮���O���s�� ��>���b�t��� '��K��������� :�L���p������5� ��Y��� ��$��H ��U~�1�� g�� 2�V� z��?�c��
/��VISBCK�������*.VD�/[/�FR:\�F/�.�Vis�ion VD file�/��/�/� ?�)?�/:?_?�/�? ?�?�?H?�?l?O�? �?7O�?[OmO(O�O O �ODO�O�OzO_�O3_ E_�Oi_�O�__._�_ R_�_�_�_o�_Ao�_ Rowoo�o*o�o�o`o��o�o�o�oO��M�R_GRP 1G���L4uC4 w B�8p	 �����|�p۬B���D��f�nӺMT� ��� ����u �y�q���r�x%��t�A�5s�s_�J�N���L1��L�5�M���H^/E��L�������p@4��B���Az�?��Bf��9�f����B��B��B
�B���B�����F@ %���-���g�fF6��D�MqD�� �BT��@���❍?@�u�Ï6���؝���5��5�����Ɵ���ß��� ��A� ?�M��r�����������  @���@�h0?�\	@�B�ɯ�����8� #�\�G���k��������ڿ���4uBH8p 9��:�L�^����̲Z��W[�a`�w���;�A@O�~��@�33@���'�\����ɿ� Ɋ��"߼�I�[�F���jߣߎ��߲�<�G��=�<�m�]<�+=~��m<c^��8e�N7��7���7�x7;�51���:���7�Tp��t2�pY�p��p��O��O��w�⮪�p �pO�0'���t���-��� C��#�1���Y���� ����������0T ?xc����� ��>)bM ��N�P�^�Z�� /�+//(/a/L/�/ p/�/�/�/�/�/?�/ '??K?X9�X?~?�? �?i��?�?=?�?�?O OBOTO;OxOcO�O�O �O�O�O�O�O__>_ )_b_M_�_q_�_�_�_ �_�_oo��7o�{� %�7��o[��o��o�_  �o$H3X~ i������� ��D�/�h�S���w� �����㏩�
���.� �R�=�v�a�s����� П����ߟ��(�N� 9�r�]���]?��̯ޯ �?�{�$�J�5�n� U���y���ȿ���׿ ���4��D�j�Uώ� yϲϝ����������� 0��T�o-o��Qo�� uo�o�߫o��o5�G� P�;�t�_����� ��������:�%�^� I���m����������  Ǐ!�ZE~ i�������  D/hS�w ������
//./ @/�d/��/s/�/�/ �/�/�/?�/?<?'? `?K?�?o?�?�?�?�? �?O�?&OOJO5OnO YOkO�Ok�}��O���O ����1_��U_�O�_ y_�_�_�_�_�_o�_ 0oo@ofoQo�ouo�o �o�o�o�o�o�o, Pq;�[�� �����:�%�^� I�[��������܏Ǐ  ���6��Z�l�~� E/O����؟ß��� ��2��V�A�z�e�w� ����ԯ������� ,�R�=�v�a������� ������O�O'�I_K� _7_9_?ϥ�o_տ�� �������8�#�\�G� ��kߤߏߴ������� ��"��F�1�j�U�g� ��g�������� �B�-�f�Q���u��� ����������, P;t�M���� ���k(L3 \�i����� ��$//H/3/l/W/ �/{/�/�/�/�/�/? �/2?D?�e?/ϩϛ? eϿ?�ϟ?��
O%?.O ORO=OvOaOsO�O�O �O�O�O�O__(_N_ 9_r_]_�_�_�_�_�_ �_��o�_8o�_\oGo �oko�o�o�o�o�o�o �o"F1C|g �������� �B��;�x�c����� ��ҏ�������>� )�b�M�_��������� ��˟���:�%�^� I���I?[?��?ٯ�? �?��?3��?Z�u�~� i�����ƿ���տ�  ��D�/�h�Sό�w� ���ϭ�����
���.� �_oo'߈�s߬ߗ� �߻������*��N� 9�r�]������ ������8�J�\�n� 5�������������� �� F1jU� y������ 0T?xc��������$FNO ������
F�0!   T�1 �D|���RM_�CHKTYP  ����������!OM _MsIN" ����N ��  X�SS�B_CFG H�� ���{/��r#�/�/�T�P_DEF_OW�  ��-"�(I�RCOM! �/�$�GENOVRD_�DOC&�ѡ<T[HRC& d5d4o_ENB�/ 0�RAVC_GRP� 1Id'�! X ��?��?�?�?�?�? O&OOJO1OnOUOgO �O�O�O�O�O�O�O"_ 	_F_X_?_|_c_�_�_ �_�_�_�_�_�_0o2�ROUp0O�Q ������"��8�?T��o3o|o��o�o��  D3A�1�ov/��@r�|B�ҡrĩoi4o�g0SMTm3Pt=��e����HOS�TC]"1QOip [��o 	�x�{��0�'�O�eC�t���������b��ۏ����4�5�Ȁ	�anonymous8�f�x�������� ���.�P�ʏ7�I� [�m���������ǯٯ ��:�L�!�3�E�W�i� ��ʟܟ���տ$��� ��/�~�@�e�wω� �Ͼ���������� +�z�����D߲ϗ�� ����������'�9� K�]�߁��ϥ���� ����<�N�`�r�t�Y� ��}������������ ��B�0��gy ������"�4�6 j�?Qcu��� �����T)/ ;/M/_/q/���� ��/,??%?7?I? �m??�?�?�?�// (/�?O!O3O�/�/�/ �/�?�O�/�O�O�O�O _Z?/_A_S_e_w_�O �?�?�_�_�_�_j}�q�ENT 1ROk� P!�_Eo  @p3opo_o�oWo�o {o�o�o�o�o6�o Z~A�e�� ��� ��D��h� +�=���a���揩� 
�͏�@�/�d�'��� K���o�������ɟ *��N��r�5���Y��k�̯��𯳯�ת?QUICC0!����p�3�1q�M�_����3�2�������!?ROUTER�����`�!PCJO�Ga�<�!19�2.168.0.�10:�gNAME� !"j!RO�BOT��nS_C�FG 1Q"i ��Aut�o-starte�d`DFTPkO HтO�_s߸O�ߩ߻� ����$_��'�9�\� J��߁������JF !�3�E��Y�{�1�b� t�����g�������� '���:L^p� �QOcOuO� O� $6HZ)~�� ���k�/ /2/ D/V/����/��/ �/�/
??��/R? d?v?�?�/�???�?�? �?OOg/y/�/1O�? �O�/�O�O�O�O�O�? _&_8_J_mOn__�_ �_�_�_�_)O;OMO_O a_Fo�Ojo|o�o�o�o �_�o�o�o/o�o�o Tfx���_�_o !o#�Wo,�>�P�b� t�C������Ώ��� ���(�:�L�^��� ���ʟ�� �� $�6��Z�l�~����� şG�د���� ����T_ERR S���.�>�PDUSI�Z  �^���U�>n�WRD �?ը��  �guest \�����ҿ���Ͽ��SCD_GROU�P 2TM� ����1�!��L9_N��  ��>R�	 i-	��v�����E E�ATSWILIB���\�N�ST �4�@��bǀ�}�FRS:�T�TP_AUTH �1U=�<!iPendan�޶�����!KAR�EL:*�(�:��KCO�_�q�G�V�ISION SE!T8��ߦ��!���� ��D�"��:�4��X��j������CTR/L VM�����
��FFF�9E3�璉��D�EFAULT-��FANUC W�eb Server-�
�Ė�����������������<�WR�_CONFIG �W�����-�>�IDL_CP�U_PCL���B�ȩ�g �BHMM�INXE�lGNR_IOG�|���S�O �NPT_SIM_�DO��TPM�ODNTOL� >�_PRTY�g�KOLNK 1XM�	�-?Qcu���MASTEҜ ���	O��O_gCFG��UO��|��CYCLE���F�_ASG 19Y*�
 �\/ n/�/�/�/�/�/�/�/��/?"?4?F?�/"N�UM{�Q�{��I�PCH/���RTRY_CNL�Q���SCRN_UP)D{�,�U� ����ZM�r�O����$J23_DS/P_EN��M���~@OBPROC$C���JOG4�1[�M� @��d8��?�Q;�OQ??>ZCPOSREDO��KANJI_�K���CM��3\*�x�E�O�ECL_Lw �l2�?�@EYLOGWGIN����|A�U��$LANG?UAGE ��g�F� �Q>�LG��2]�ﱢ����xRBа���Pm ����'0�H���0��MC:\RSCH�\00\.��PN_DISP ^M�॔��|�z�<�LOC��^Dz�=#��{�iPBOOK  a�>'}@���������`XJi�o�o�o�1~D}7xVy�	�e�i��Me��}b�G_BUFF 1-`�2��� �b�����'�T�K� ]�����������ɏ�� ����#�P�G�Y����)d`@DCS b>�m =���S|�������� �8C��I�O 1c:+ 	O]����]�m���� ����ǯٯ����!� 5�E�W�i�}�������@ſտ����8�E� _TM  9kdC� Y�k�}Ϗϡϳ����� ������1�C�U�g� yߋߝ߯����߾t=��SEV�09m7�TYPC�U�6�H�Z��}�ARS| R_�s�2�FL 1dF��0�Ο��������(�L:�k�TPfPC�%�}rmNGNAM$D�e	��UPS1`G�I�5 Q�5��_L�OADA@G %�9j%CAL_T�C���D
MAXUALRMl7�z8 ����3�0�Tq C4ae��i�~S tb@g@f:+ �w	%�����- Q<uXj�� ���/�)//M/ 0/B/�/n/�/�/�/�/ �/?�/%???[?F? ?j?�?�?�?�?�?�? �?�?3OOWOBO{O�O pO�O�O�O�O�O_�O /__S_e_H_�_t_�_ �_�_�_�_o�_+o=o  oaoLo�ohozo�o�o �o�o�o9$]�D_LDXDI�SA��E�6�MEM�O_AP��E ?=��
 �fy ������&�8�~ ISC 1g�� �P��Lt���� ��O؏Ï��� �2� ��A��z�e������� ԟU�㟷��.��R� 9�v�������k�Я�� ��ۯ�*���9��r� ]�������̿M�ۿ�� �&��J�1�n��}� ��c��ϳ������"� ��1��j�Uߎߠ�Y��_MSTR h��ݳ�SCD 1i�}�����&��J� 5�n�Y�k������ ������� �F�1�j� U���y����������� ��0T?xc ������� >);t_�� �����//:/ %/^/I/�/m/�/�/�/ �/�/ ?�/$??H?3? X?~?i?�?�?�?�?�?��?O��MKCFG� j��O��L_TARM_5Bk��wKB C��p�NxpMETPU܅pB����NDSP_CMNT�EpI@CF�E�� l�ނ�NBKA_T�EP�OSCF�G�NP�RPM�O�HPST�OL 1mc�4@@<#�
�Q	A�U �_�W�_�_�_�_o�_ �_<oo0oroTofo�o �o�o�o�o�o�a�A�SING_CHK�  \_$MODAQhCn;O�GKJNu�DEV 	��	�MC:~|HSI�ZE�@���NuTA�SK %��%$�12345678�9 ��uLwTRIoG 1o�� �F3%��OL�  1�r�U����vYP�q]����MsEM_INF� 1poG �`)AT&�FV0E0���)�ށE0V1&A�3&B1&D2&�S0&C1S0=>�)ATZ��J�1�HN�v��j���-�A��Ο���ٟ�(� ܏M� ��$�6��� Z�˯�����%�� I�[�B��2�D���h� z������¯3�j�W� ����HϱϘ����� ��߾�п���e�� ���Ϛ߿�r��ߞ�� � �=����s�&�8� J߻������(���� ��K��o�V�����X� ��|����#��G Y��}0��\�����#NONITO�R�@G ?�{  � 	EXEC�1C>2D3D4�D5D�F7D8
D9C?��C �O�[�g�s ���������2�2�2�2��2�2�2�2�(2(2(3�3�3ONqR_GRP_SV 1qˉ�,�(q>�9�?��h���?���<��@�g,Ѯy}�q_D���~0APL_NAM�E !�E;0��!Defaul�t Person�ality (f�rom FD) �-DRR2�! 1r�)deX)dh�;1�AX dO�?�? �?�?�?�?OO%O7O IO[OmOO�O�O�O�O�O�O�O	X2�?-_?_ Q_c_u_�_�_�_�_�_=r<_�_oo/oAo Soeowo�o�o�o�o}x�R�" 1w39jp=\@r0 ���@r��a @D�  &q?�s�a?@pq�@qAI�Ez � 3qqEw;�	l~'r	 0Ap�er@es_qp�{t��{t� Ki�K��J���J����J�4�J~���Ezvq�^q�P���|�p@�z��r�f�@�S���/q��s�=�N���
������T;f�
�����p�*  �_p  �U�>Q���U���?��?�����OO�����R�����(q����Buʍ�|}  ����pj  T�������܏ 	�'� � C��I� �  {��ߍ:�Èg�?È=�����r@�����~q��D*�rÈ��~N_0�  ''��q(��@a�@�t�E@4�@8���pCP�KCa�fa�\�B`��Cd�p�@�V��voo$~�}����wAAV���_0ϡ*��pp�qD8u�����5� �Y��}�� ��t O� �ru �4 ������Ӄ� �::u�qp�p �?�ff Q��Ŀֿh� ������q�4�B�>������yPplϖ���xvqevم�>L������r<	�I<�g�<#�
<2���<D��<���
����s��s_��?fff?榐?&��t@T���/�?�`?U?ȩ?X�?��� ���(tk�ts�w�� �[t���߲������ ��3��W�i�T���\�F_0|���x����d������A���G�@ G��F���� t������������� +�z��O�  ڏ��(��d' 9K��`r��P����Ϣ�$ ��&/w�M/�q/\,�w��z/�/�/�/�)�2V��$-�pB�a�01?m��"�� �!71�@I�;M`B�@��@`�9�@y��?�h�? �@�3��[N��N�N�E��<�/k?�}0�>��ڟ��A�p�C�F�@�S��?u�X������@�t��%�h�?�K�G��Gk�nF&�Fצ�pE,8{�? �F�ZG����F�nE�D�E,ڏO@����G��F7���F��ED�� _��/tO_O�O�O�O�O �O�O�O__:_%_J_ p_[_�__�_�_�_�_  o�_�_6o!oZoEo~o io�o�o�o�o�o�o�o  D/hSe� �����
��� @�+�d�O���s����� Џ��͏��*��N� 9�r�]�������̟�� �۟���8�#�5�n��Y���}�����گŮ(��13�jiꯣ��y��ӥ3Ա��<��4 ��7�I���P�c�u�W��jb����1w�����������@���C�1̤P��	PuΔ����� ������#�М��� >�)�A�M�_�5$x�B� �߮��������ņ ��{�5�C�U�y_�q� �������e����-��Q�?�u�_�2v�0�$��G��ߢ� B !!� B
�CH � K���� &8J���~@������$��E� � �ў�c�%
 �0BT fx��������//�:
 ���o�x}��$M�SKCFMAP � ���� ��
��-S#ONREL  g��j!��S"EXC/FENB�'
h#�%ε!FNC�/�$JO�GOVLIM�'dt� �"dS"KEY�'u5S"RUN�,�5S"SFSP�DTY���&�%�#S�IGN�/�$T1M�OT�/�!S"_C�E_GRP 1x��j#\ϯ�?ǯ OOe�??O�?cOO XO�OPO�OtO�O�O�O _)_�OM__q_�_:_ �_^_�_�_�_oo�_ 7o�_[omoTo�o^S �TCOM_CFG 1y`-�o�o��o
�a_ARC_�"g��)UAP_�CPL�$NOCHECK ?`+ f�lxj| ����������0�B�T�f�x��+N�O_WAIT_L�w7f%�2NT�az�`+ʁ_ERRr�2{`)��� �o#�5�G�S�9#k�}�^ItT_MO��|��, nr�oȟ��_PARAM�2}`+�	���~g���E� =��345678901_�q��� Z������������د0 �2��}g�d�v��	���JsUM_RSPACE]/ӿݴ��$ODRDSP�sz6�(OFFSE?T_CART9��DIS��PEN_FILE<�z1�a���pOPTION�_IO?�PWO_RK ~�7�# �Э�t��
g�8������	 ������t����RG_D?SBL  ��#�6��RIEN�TTO� ��C��i!=#�p�UT�_SIM_D{��g":"�V��LCT ԍ�����a��>��_PEXE=���RAT���&�%M0��>�UP ������%�7��[�i���$�2�3r)d�eX)dh���X d�������� ����
��.�@�R�d� v���������������$2��HZl ~��������<7&8J\n �������'���0O�1w(��O�(�_Ҙ��20 �Ԧ  � @D�  .!?��4#!?��6!��D4  EzP#Ijd,�;�	lF"	 '0��"@�#~!�* ��$��$1�H)�!H,�H�8�Hm�G�?	{G�8�$�g��~f��/ <1�C�Z�1�Z�� 3N!-?���*  �p � �L0>H0� # �+=C?U2�]��-�B]�Btr�«{���¼�2?�?�2G!�31�])�a/1�@�  �@��j  K0�&F��DO~e	'� � bB�I� �  ����==���8�O�K`�@�O�@ �>��OIK�0�N�&ykN ._4Q'~�HT,1o0CZ�fZ�S0BW0*>S_eR\�IJ�a��@uA�&o�o$�-���{gAu@�Z5P�QIJ �AeJ" W%3O0ooTo?oxocm��� �t �O� ru �4 ��b<�e��� :�5�����0 �?�fAf�qk�o�o�o�ʈ3��Q8��Saz>��`�agiP����g�Q�!�&�5�>L��@�32<	�I<�g�<f�<2���<D��<��`���/�5"��|~r`?fff?�@�?&<�kd@T��N�?�`?U��?X�^���R 7�G$fi6%��4'�� � z$�я
���.�� R�=�v���s������� �͟�}�������`�~��G�@ G�0 ��������ί���� �(��L�7��Rn�1� _��?��?#��G�� ��4�F�X�j�	�ϑπ+��ϯ���������R�4��TEߖ��l�xߐ�{�?�ؙ�P���������uD�C��1��P'�&�1�ظ���в�V�@I��Z�M`B@���@`�9@y���?�h:� ��@�3�[N���N�N�E��<��/����>���ڟ�A�p��C�F@�S����8�X������@�t��%��h�°�1G���GknF&��FצpE,8�{� F�Z�G���F�n�E�DE,ڏ�*�<��G���F7��F��ED��~v�ߓ�~� ������������5  YDi�z�� ����
U @yd����� ��//?/*/c/N/ �/r/�/�/�/�/�/? �/)??9?_?J?�?n? �?�?�?�?�?�?�?%O OIO4OmOXO�O|O�O �O�O�O�O_�O3__ W_B_T_�_x_�_�_�_��_�_�^(��3�j�i	o�q��:e�U3�Ա�*o<o�q4 ��Voho�q�Pqło�ovbjb�o��o1w������m�i>,b�P|õP�rP�~�� ���o��o��Bi#���$�]�H�`�l� ~�Tԗ�aߏ͏�� '�=i�u������T�b�t�y~���Ɵ��ʟ؟ ꟬r���2�L�:�p�h^���~z2��$�f'G����`B?�3��B)�CH4��`j� ��+�=�O�a�s�ɳ��������ӿ���*�d��`�`��r�����e
 �� O�a�sυϗϩϻ��� ������'�9߸�)�� ����x}���$PARAM_MENU ?���  �DEFPU�LSEE�	WAITTMOUT���RCV�� �SHELL_WR�K.$CUR_S�TYL����OsPT���PTB���C��R_DECSN�ЅuX�R�d�v� �������������/�*�<�N�w�r�US�E_PROG �%��%s�����CC�R���u����_H�OST !��!����T�p��)���+e��_T�IME��1��  �r�GDEBUG�/ �ۇ�GINP_�FLMSK��	T�R��PGA�  2����CH���TYPE~��� r�l������� � //;/6/H/Z/�/ ~/�/�/�/�/�/�/? ? ?2?[?V?h?z?�? �?�?�?�?�?�?
O3O��WORD ?	>	RS� �S/PNS�U��oBsJO��RTEL �0TRACECToL 1����� �p ��p�p�N�FDT� Q���@�@�D(���P�R6��smU�q-P )�3R%�WP0RP8R�P@RP�R�R�	T	T		T	T*	T	T	T	T1 �R	T	T	T�	T	T	T	T�	T	T=�R	T�	T�R!	T"	T#�	T��R&	T''� E_W_i_{_�_�_�_�_��_�_�_oo/o	T%TIhQ(	T)	T*	TU+	T,	T-	T.	T/	T0Qocouo�o�o �o�o�o�o�o) ;M_q���rQU1	T2	T4	T5	TU6	T7	T9	T:	TU;	T<	T=	T>	T%?	T@	TY�� ����!�3�E�W� i�{�������ÏՏ� ����/�A�S�e�Q ]Q�c�u��������� Ͽ����)�;�M� _�qσϕϧϹ����� ����%�7�I�[�m� ߑߣߵ��������� �!�3�E�W�i�{�� ������������� /�A�S�e�w������� ��������+= Oas����� ��'9K] oE������� �/#/5/G/Y/k/}/ �/�/�/�/�/�/�/? ?1?C?U?g?y?�?�? �?�?�?�?�?	OO-O ?OQOcOuO�O�O�O�O �O�O�O__)_;_M_ __q_�_�_�_�_�_�_ �_oo%o7oIo[omo o�o�o�o�o�o�o�o !3EWi{� �������� /�A�S�e�w������� ��я�����+�=� O�a�s���������͟ ߟ���'�9�K�]� o���������ɯۯ� ���#�5�G�Y�k�}� ������ſ׿���� �1�C�U�g�yϋϝ� ����������	��-� ?�Q�c�u߇ߙ߽߫�����������$PG�TRACELEN�  ��  �_������_UP �����@�H�,��A��_CFG M�@�*���A��m�#� m����m�U�DEFSPD� �`��q#����INX�TRLW �`���8}����IPE_CON�FI\��@���@�m���LI�DY�`�<�GR�P 1��*�����@�
=�[����A?C�C�
�XC)��Bg����#�����d}����/�/�� 	 ��������� ´����B  8N8r���> �6>7��D���� ='?�=)��� �O:s^���~���  Dz#/��
/G/� W/}/h/�/�/�/�/�/ �/?�/
?C?.?g?R?��?��
V7.1�0beta1m���0B=q�2`�ff@��2>�{���1=����1�A>ff�1@�f�f�2�\)�2D�_�?�  A@	AL�0�1Ap�3�ș?`7OIO[OmO|K�����,��?�O|?�O�O _ _9_$_6_o_Z_�_ ~_�_�_�_�_�_o�_ 5o oYoDo}oho�o�o �o�o�o�o&/1�o U@R�v��� ����-��Q�<��u����?�3F@  ��������@��M� �0�&�N�`��O�O�O ������ޟɟ��&� �J�5�G���k����� ȯ���ׯ�"��F� 1�j�U���y������� ���ͿB�-�f� Q�cϜχ��ϫ����� ���,�>�)�bߍ��� я�߭������� A�:�e�w�������C� ������������6� !�Z�E�W���{����� �������� 2V Aze������ �
�.R=v as������ //</N/yߋ߽߇/ �/���߻/�/�/-�&? Q�c�u��?//�?�? �?�?�?�?�?"OOFO 1OjOUOgO�O�O�O�O �O�O_�O0_B_-_f_ Q_�_u_�_�_��_�_ �_oo>o)oboMo�o qo�o�o�o�o�o�o (S/e/w/�/s�/�/ �/?�? ��=?O? a?s?l���{����� ؏�Տ���2��V� A�z�e�w�����ԟ�� �����@�R�=�v� a����_��Я���� �*��N�9�r�]��� ����̿���ۿ�? Qc�_ϙ���� �������)�;�M�� X��|�gߠߋ��߯� �������	�B�-�f� Q��u��������� ���,��P�b�M��� ������k����� :%^I�m� ���� +�=�O� 9K�ϗϩϟ��� ���'�9�2/�// h/S/�/w/�/�/�/�/ �/
?�/.??R?=?v? a?�?�?�?�?�?�?�? OO<O'O`OrO���O �OWO�O�O�O�O_&_ _J_5_n_Y_�_}_�_ �_�_�_)[%o7o�q���o�o��$�PLID_KNO�W_M  ����Q�dSoV ���`��O! 3�_WBT��R-��cM_GRP 1���j& dzp��oo$tv�t_���d��d M`�z	�}{�v,�S��e �o�C�?���c���ۏ �������5��h�e� )�K���u��������� ���+���g�;���`I�[���Ӯ�aMR�sŎ�}T�Uxa|O  xb3�E�Y�T�*���N� `�r��������̿.� @�U�P�&ψ�J�\�n� ���ϼ϶���*�<�Q�`L�"߄�F��ST�q�1 1�����v�`0� @��� �U�������H�+�=� ~�a�s�������� �����'�h�K�]������2�����Q�<����3����������4/A��A5Zl~���6������7�
.��8GYk}�ӿMAD  $��� ��PARNU/M  ��|����SCH� �
�<'!J)�c\%UPD�/%�q�/�$��_C�MP_�p�m`�'��e�$ER_CHK�%���j�"�/��+RS��o�a_M�O�.?@5_*?�__RES_G�А�� */���?�?�?�?O �?%OO*O[ONOOrO@�O�O�O{7���<�? �O}5
 �O__3Y  &_E_J_3� e_�_�_ 3� �_�_�_3F�_ oo3�"oAoFo2�V 1��e�q"@�cX��`P�`�`W���`l�` @cV���`�@2THR_�INR���rr5d��fMASS�o Z��gMN�osMON�_QUEUE Q��u�&�p��p�N� U1N v�+cp�ENDeqg?yEX1E�u� BE�po>`sOPTIOlwp;�cpPROGRAM7 %Cz%bp�o�+/arTASK_I���~OCFG �C/7�j�DATuA���s�@��2�������'�я J�\�n���+�����ȟxڟ쟟�INFO������Rt��@�R�d� v���������Я��� ��*�<�N�`�r���Ж�������� ��Ii�� DIT �s�ϛ�WERF�L�x�c��RGAD�J ���A�  ]�?v�i��aA�cq�n����'�?���v�<��/�%���5ȲO��±��2���!�t 	 h���b�����Ard�t$B�v��*U�/W� **�:`�P�bր�;����ҍ՝߉5��NӼ� ���ߕ��������� ��A�7�I�[���� �������=�����v� !�3���W�i�{����� ��������o� ASЇ�� � �C�'I��U�y��RIORITY� w�&�E�MPDSP�q3ϱUw-��;OG�_TG0�W��Gz�TOEp1���� (!AF��`Ef09/D'!�tcpD/l-!�ud[/�.!iccm�/�o�XY��������)� 0m��/
?����/3? 5"?_?F?�?j?|?�? �?�?�?OO�?7OO�[OmO*D�PORTT�q���%E��_CARTREP��p���aSKSTA�x�zSSAV?p����	2500H809�(����D������`.�kY_xk_i�PURGE�p�B0��yWF�PDOU���W2 �T��J�WRUP_DEL�AY ����TR_HOT��b��8o��UR_NORMA�L�(o}oLfSEM�I[o�o�oqQSK�IP���� x kg);M} ~l������ � �2�D�
�h�V��� ����v����ԏ
�� .��R�@�b������� r�П������ޟ(��N�<�r�������$�RBTIF���R�CVTM�$����DCRƳ��l��qB
�B}��>A��@��_��"���x��$��Q�V����HU���o���6�`�\ �<	�I<g��<#�
<2���<D��<���
r�Y�¿Կ  ֿ��� �2�D�V� h�zόϞϰ��ϭ��� ��
����@�+�d�G� �ߚ�ݿ��������� �*�<�N�`�r��� �ߺ���������� 8��\�n��ߒ����� ��������"4F XC�U��y��� ���0B��f x������� //,/P/;/M/�/ q/�/�/�/�/�/?G Y:?L?^?p?�?�?�? �?�?�?�? O�/$OO HO3OEO~OiO�O�O�O �O?�O_ _2_D_V_ h_z_�_�_�_�_�_�O �_�_oo@o+o=ovo Yo�o�o�O�o�o�o *<N`r�� ��o������ 8�J�-�n����o���� ȏڏ����"�4�F��X�j�y��GN_A�TC 1��� �AT&FV�0E0y�AT�DP/6/9/2{/9��ATAy��,AT%G�1%B960���+++ޟ,ّH��,�IO_TY�PE  \�ƣ�e�{�REFPOS�1 1�G� O x�f���_� Ư[���������B� -�f����%���I���俒�����ҿ3�� W��{�ϟ�:Ϝ��� p��ϔ�߸�A�����  �:ߛ߆߿�Z���~� ���=���a��߅�  ��D�V�h����� '���K���o�
�l��� @���d��������� ��
kV�*�N �r��1�U �y&8r�� ��/�?/�</u/ /�/4/�/X/�/|/�/ �/�/;?&?_?�/�?? �?B?�?�?x?O�?%O �?IO�?�?OBO�O�O �ObO�O�O_�O_E_ �Oi__�_(_�_L_^_ p_�_o�_/o�_So�_ wooto�oHo�olo�o �o�o�o�os^ �2�V�z�� �9��]����g�y�2 1���.�@�z� ����"�@�ۏd��� a���5���Y��}�� ����ş��`�K���� ��C�̯g�ɯ���&� ��J��n�	��-�g� ȿ��쿇�ϫ�4�Ͽ 1�j�ώ�)ϲ�M��� qσϕ���0��T��� x�ߜ�7ߙ���m��� ����>�������7� ����W���{���� �:���^������� A�S�e��� ��$�� H��li�=� a����� hS�'�K�o �
/�./�R/�v/ /#/5/o/�/�/�/�/ ?�/<?�/9?r??�? 1?�?U?�?y?�?�?�? 8O#O\O�?�OO�O?O �O�OuO�O�O"_�OF_ �O�O_?_�_�_�___ �_�_o�_	oBo�_fo�o�o%o�o����3 1���[omo�o% IOom�,�� b����3��� �,���x���L�Տp� ������/�ʏS��w� ���6�H�Z������� ���=�؟a���^��� 2���V�߯z������ ¯��]�H������@� ɿd�ƿ����#Ͼ�G� �k���*�d��ϰ� �τ�ߨ�1���.�g� ߋ�&߯�J���n߀� ����-��Q���u�� ��4����j����� ��;�������4����� ��T���x�����7 ��[���>P b���!�E� if�:�^� �/���/e/P/ �/$/�/H/�/l/�/? �/+?�/O?�/s?? ? 2?l?�?�?�?�?O�? 9O�?6OoO
O�O.O�O�RO�O�o�d4 1� �o�O�O�OR_=_v_|O �_5_�_Y_�_�_�_o �_<o�_`o�_ooYo �o�o�oyo�o&�o #\�o��?� cu��"��F�� j����)���ď_�� �����0�ˏݏ�)� ��u���I�ҟm����� �,�ǟP��t���� 3�E�W����ݯ��� :�կ^���[���/��� S�ܿw� ϛ������� Z�E�~�Ϣ�=���a� ���ϗ� ߻�D���h� ��'�a��߭��߁� 
��.���+�d��߈� #��G���k�}���� *��N���r����1� ����g�������8 ������1�}�Q �u���4�X �|�;M_� ��/�B/�f// c/�/7/�/[/�//?<�O T5 1�_�/ �/??j?�?�/�?b? �?�?�?!O�?EO�?iO O�O(O:OLO�O�O�O _�O/_�OS_�OP_�_ $_�_H_�_l_�_�_�_ �_�_Oo:osoo�o2o �oVo�o�o�o�o9 �o]�o
V�� �v��#�� �Y� �}����<�ŏ`�r� �����
�C�ޏg�� ��&�����\�埀�	� ��-�ȟڟ�&���r� ��F�ϯj�󯎯�)� įM��q����0�B� T����ڿϮ�7�ҿ [���Xϑ�,ϵ�P��� t��ϘϪϼ���W�B� {�ߟ�:���^����� ����A���e� �� $�^�����~���� +���(�a���� ��� D���h�z�����' K��o
�.�� d���5?-46 1�8?��. ������/� /N/�r//�/1/�/ U/g/y/�/?�/8?�/ \?�/�??}?�?Q?�? u?�?�?"O�?�?�?O |OgO�O;O�O_O�O�O �O_�OB_�Of__�_ %_7_I_�_�_�_o�_ ,o�_Po�_Mo�o!o�o Eo�oio�o�o�o�o�o L7p�/�S �����6��Z� ���S�����؏s� ���� ����V��z� ���9�]�o����� ��@�۟d�����#� ����Y��}����*� ůׯ�#���o���C� ̿g�𿋿�&���J� �n�	ϒ�-�?�Qϋ� ����߫�4���X��� Uߎ�)߲�M���q��� �ߧ߹���T�?�x�� ��7���[���������>���b�HZ7 1�e�!�[����� ���!��E��B{ �:�^��� ��A,e �$ �H��~/�+/ �O/��/H/�/�/ �/h/�/�/?�/?K? �/o?
?�?.?�?R?d? v?�?O�?5O�?YO�? }OOzO�ONO�OrO�O �O_�O�O�O_y_d_ �_8_�_\_�_�_�_o �_?o�_co�_�o"o4o Fo�o�o�o�o)�o M�oJ��B� f�����I�4� m����,���P���� �����3�ΏW��� �P�����՟p����� ����S��w���� 6���Z�l�~����� =�دa����� ����� V�߿z�Ϟ�'�¿Կ � ρ�lϥ�@���d� �ψ���#߾�G���k��ߏ�u���8 1� ��<�N߈����*�0� N���r��o��C��� g������������ n�Y���-���Q���u� ����4��X��| );u���� �B�?x� 7�[���� >/)/b/��/!/�/E/ �/�/{/?�/(?�/L? �/�/?E?�?�?�?e? �?�?O�?OHO�?lO O�O+O�OOOaOsO�O _�O2_�OV_�Oz__ w_�_K_�_o_�_�_o �_�_�_ovoao�o5o �oYo�o}o�o�o< �o`�o�1C} ����&��J�� G������?�ȏc�� �������F�1�j�� ��)���M���蟃�� ��0�˟T����M� ����үm�������� �P��t����3�����ߴ�MASK 1����� ���?XNO  ��~�MOTE  /�����e�_CFG ��lͷ���PL_RANGh�b�p��POWER �����x�SM_D�RYPRG %�l�%i����TAR�T ����UME_PRO�� �{����_EXEC_E_NB  `�tɏGSPDTЖО����TDB����R�M����MT_�T���j��OBOT�_NAME �l�j�׹OB_O�RD_NUM ?����=�H809  `����	d�H	��\췰���� ,��:��	@���D|����PC_TIMoEOUT�� x�oS232��1�0���� LTE�ACH PEND�AN������)��[�R� M�aintenance Consb��&�_�"B�T�KOCL/C.Д�r��5��� No Use��r���]���NPO������v���CH_�LW��lβ�	�a0MAVAIL�w�����t���PACE1 2�l� +���	������p�8�?��,	;, q�i���� �	�-OA/b/%/ ��/)0�4��-�� �	/{/-/O/A?b?%?@�/�??�?:�2���/�/?�?+?M? \O}O@O�O�O�O�O�;3�?�? OO$O�OHO jOy_�_]_�_�_�_�_�;4�O__/_A_�_ e_�_�o�ozo�o�o�o�;5o(o:oLo^o �o�o����
����;63EWi {)���Џ񏴏�'��<��;7P�b�t� ����F���ޏ��џ #�D�+�Y��;8m�� ������c�ٟ��
�+���@�a�H�v��;h �Nl� m��
Ӱ ¿����� %�7�I�[Ϲ(˧~ͱ� ����S����d��ؿ ��*�<�N�`�r߄� zόϞη/�ߓ����� �0�B�T�f�x��� �߼���������� "�P�b�t������������������
� `n� @�S�� a=�E��!*� ����
��)G �/q�MWi� �����7/I/g/ /O/�/�/m/w/�/�/��/�/��
�R?�;_MODE  ��^h9S ���A?����ޯ}�?�?J�	OAO�DCWOR�K_ADx=	5���AR  ��𚠏@FOy@_INT�VALx0����:R_OPTION�F� �5`V_D�ATA_GRP �2�����D9�P .O_*O>_)Y+?k_Y_ �_}_�_�_�_�_�_�_ �_1ooUoCoyogo�o �o�o�o�o�o�o	 ?-OQc��� ������;�)� _�M���q��������� ˏ��%��I�7�m� [�}�����ǟ���ٟ ����!�3�i�W��� {�����կï�����/�1�$SCAN�_TIMw1I��5�I�R �(�3�0(�L8�ѰѲ�34Q	���1���:�3_�����?��Ӳ2Ĉ���d����/R�� @���Q�c�u�RU0�D� �P��0[ � 8�@��������D�����+�=�O� a�s߅ߗߩ߻��ߒ��1B����#����S����;��oRT���1p���?t��DiD��>��  � lӲ�1 �񘱐����������� ���#�5�G�Y�k�}� �������������� 1<��Sew� ������ +=Oas��� ���>P�� /2/ D/V/h/z/�/�/�/�/ �/�/�/
??.?@?R?�d?v?�?�?�5�?  0�2'���?�?O#O 5OGOYOkO}O�O�O�O �O�O�O�O__1_C_ U_g_��_�_�_�_�_ �_�_	oo-o?oQoco uo�o�o�o�o�o�o�o v_�_/\n� �������� "�4�F�X�j�|�����`��ď֏�7�?  � 
��.�@�R�d�n��� ������ɟ۟�����#�5�G�Y�k�}��� 葯�è�ί�� ��(�:�L�^�p����ɶ����¿������ ����	�12345678����������02�D�V�h�z��������������� ��0�B�T�f߭��� �߮����������� ,�>�P��t���� ����������(�:� i�^�p����������� ���� A�6HZ l~������ �+ 2DVhz ������
/ /./@/R/d/v/�/�/ �/�/��/�/??*? <?N?`?r?�?�?�?�����?�?�3�/OO�)OMyCz  B}p��   �Qx�2���:�$SCR�_GRP 1�(��e@(�l��0�@} � ۱��	 �C�A�B�D�1����I���F�O�O$_I}[���C�PP�������fX![w\L�R Mate 2�00iC �90���U�LR2CA ���C���
�X��S�AշV�wS��!Q�J�Ai	�RLo^opo�o�o�lް��@5n߲�o �O!_
�G�?���@`�o�=Hv?Fh�-,�IB�K@���r��t�AA\@�  @����A@WP�  ?~�6��rHK@G��z��AF@ F�` q�y�p��������я �����?��}�>�`j�U�g�y���B��� .�ߟʟ��'��$� ]�H���l�����ɯX^�ū��_�����e
��Y��6�@��=�ò"`��G"���B�6���90��>G��@EL_DEFA�ULT  �d�_�/�ޱ�MIPOWERFL  �E��ݲ�oWFDO� ����AERVENT �1����`����0L!DUM_�EIP��p��j!AF_INE�<���!FTdϽ������!�o� ����-�!RPC�_MAIN.�غ8�y�@�VISI��y�h���!TP�ГPU��w�d���!�
PMON_PR'OXY�z�e �]����+�s�fL��!RDM_SRV��rw�g����!RҸd�|�h��A�!
B��Mt�t�i0���!?RLSYNC�����8|���!ROSc� �4��%�� I��(r�^� ����'�  o6HZ������/�5/;�ICE_KL ?%K�� (%SVCPRG1:/�*l%lCD�/�-3�/�/q 4�/D�/q 5�/�/q 6"?'?q 7J?O?q �T�?�,9�?�;n$��? q!t/�?q!�/Oq!�/ ?Oq!�/gOq!?�Oq! <?�Oq!d?�Oq!�?_ q!�?/_�!�?W_�!O _�!-O�_�!UO�_�! }O�_�!�Oo�!�OGo �!�Ooo�!_�o�!E_ �o�!m_?/Q"q X/j  
OIASwb�� �������=� (�a�L���p������� ߏʏ��'��K�6� o���l�����ɟ��� ؟���#�G�2�k�V� ��z�����ׯ�ԯ� ��1��U�@�y�d���𯿚�ӿE*_DEV� K��M{C:۸̪f�OUT������?REC 1�,u��6� � 	� �Z�  
�j�m�w_Ìϝ���Q�bĽ��������w
 �Z�6 s��_�����@�Q��+vM���Y�鰕)�{�U*��B>����������ARߋ�+�,uж��r
ت���  UxR������z�K 鰝��a鰩���d�X���n�Ȋ�?nК��7�ߌU���R��R��R��E� �&� R鰟�a�=�[鰩���`�T���n�̊�*n�u����J�e��Hc�m��k� �  ���T���ե�z��.�Tp��n���6n�1zV�����~Kܽ�*i�(�t鰞�%���Q�QZ�� U�k���R�C���q;��~N@���e�a�*�P�Q>�Ɇ
D�鰱o��N���"��iR�b鰖R��RR������5/�|�� ��!UE���nм�$n�P�����*f�hR��Q��I͂*��J��_�沕C���nйB���/?/����I���P���f�./�Q<�Q�+�&$$�/,�/R/���&��`�m�R�W鰿T�/#���R�)[6?d��n����"^?�?������=�9 �?�?�?�?"OO2OXO :OhOjO|O�O�O�O�O �O_�O0__T_B_d_ f_x_�_�_�_�_�_o �_,ooPoboDo�oto �o�o�o�o�o�o�o :(^L�p�� ����� �6�$� Z�l�N���~�����؏ Ə����2� �B�h� V���z������ԟ�
���.��>�d�<�V� 1�I̜ �?����Eѡ�   -�~জ8��_T�YPE(��FZN_CFG �^������G_RP 2���/ ,BY�AY��_D;� Bq�A��B4�RB2�} �HELL�i������ ��<���%RSU1� Ͽ���>�)�b�M� ��qϪϕϧ�����߰��(�:�I��{ ���%I�w߉ߥry`%���%% ޤ7�_��d�ߏ�~�HKw 1Ō� �� =�8�J�\����� ����������"�4��]�X�j�|�x�OMM� ƌ���}�FTOV_EN��������HOW_REG�_UI��|�IMW�AIT��-0��O�UT��	TI�M��XVA�L-_UNIT�����MON_ALIAS ?e��? ( he��� �
.�6�[m �<����� �!/3/E/W/i//�/ �/�/�/�/�/�/?? /?�/@?e?w?�?�?F? �?�?�?�?O�?+O=O OOaOsOO�O�O�O�O �O�O__'_9_�O]_ o_�_�_�_P_�_�_�_ �_o�_5oGoYoko}o (o�o�o�o�o�o�o 1C�ogy�� �Z���	��� ?�Q�c�u���2����� ϏᏌ���)�;�M� ��q���������d�ݟ ���%�ПI�[�m� �*�����ǯٯ믖� �!�3�E�W��{��� ����ÿn������ /�ڿS�e�wω�4ϭ� �������Ϡ��+�=� O�a�߅ߗߩ߻��� x�����'���8�]� o���>�������� ���#�5�G�Y�k�� �������������� 1��Ugy���H����	���$SMON_DE�FPRO ����2� *SYST�EM*  �l��"RECALL� ?}2 ( ��}tpcon�n 0 >lap�top-3jv2�48ms:139�60 ver =�>3722444�8:878185= �61 1���  }7cop�y virt:\�output\c�alptcp.pc md: o� ��</N/�5� _1/�(/�/�/�/�#rxy�//�/H@?R?�)6�/2z?��)?�?�?_?�/\toest_	0ls�?  ?�?COUO�6A�2@Etp�?~DO/O�O�Oe?�OzO��O<_N_�=?rJz�O{V_ �$4_�_�_�49�O _dvO]�_=oOo�<ErEg�]zjo�38�o�o�o }8�_d@	_��o<N�=Crl _zy�$����?  /���G�Y�l/~/ ��&+���Ώa�s���2������>�P���_��0���ӟfO xc�������$��G��Y�l�;r�frs:�orderfil�.dat�ttmp?back\={��.���ѯd�2rDb:*.*�������ޯ�H�Z��w� �emp��172.23.�254.7:17884 (���˿ݿ;}-r�*.d����࠿��C�U�h�
xy?zrate 4`��@�!�3�����i�r� �ϥ��ϣϵ�F�X��Y�frh:\sup�port\��|�=�>4148428_8:936�� ,� ����b�􏆏�ݨ�9�@K�]��dw� ��� +�����a�/��ﰴ�E�W�j�3xr�: ���|���'�����.�� }4r�az���  է�8J\o��
� %�^������ �FXk�����3 ����z��B/ T/gy�//�/�/ ���/�/>?P?c u/�+?�?�?�� �?/�?:OLO�?q/�/ ?'O�O�O�O�/�O?�O�OH_Z_k`�$S�NPX_ASG �1����}Q�� P+P�'%R[1]g@1.7o�Z?�hc%�_�_�_�_�_�_.o o8odoGo�oko}o�o �o�o�o�o�oN 1X�g���� ����8��-�n� Q�x�����ȏ������ ��4��X�;�M��� q���ğ���˟ݟ� �(�T�7�x�[�m��� �����ǯ����>� !�H�t�W���{���ο ��ؿ��(���^� A�hϔ�wϸϛϭ��� ����$��H�+�=�~� a߈ߴߗ��߻���� ���D�'�h�K�]�� ������������.� �8�d�G���k�}��� ����������N 1X�g���� ���8-n Qx������ �/4//X/;/M/�/ q/�/�/�/�/�/�/? ?(?T?7?x?[?m?�? �?�?�?�?O�?�?>O�!OHOtOWDpTPAR�AM �}U��Q �	�xJP��D�@hXOFT�_KB_CFG � �C�U�DPIN_SIM  }[��F_'_9_�@pPR�VQSTP_DS�B�N�Bu_�H�@S�R �[� &�  AL_TC�E�_�D�FTOP�_ON_ERR � �D�I�QPT�N U`�A�RRINGo_PRM�_ �@�VDT_GRP �1ʝI�P  	 �G�HZolo~o�o�o�o �o�o�o�o# 2D Vhz����� ��
��.�@�R�d� v���������Џ�� ��*�<�N�u�r��� ������̟ޟ��� ;�8�J�\�n������� ��ȯگ����"�4� F�X�j�|�����ǿĿ ֿ�����0�B�T� fύϊϜϮ������� ����,�S�P�b�t� �ߘߪ߼�������� �(�:�L�^�p��� ��������� ��$� 6�H�Z�l�~������� �������� 2D khz��������
1.�CVP�RG_COUNT��F�a�E\EN�B'oWM��D�_�UPD 1�[8  
E�B�� �%/ /2/D/m/h/z/ �/�/�/�/�/�/�/
? ?E?@?R?d?�?�?�? �?�?�?�?�?OO*O <OeO`OrO�O�O�O�O �O�O�O__=_8_J_ \_�_�_�_�_�_�_�_ �_oo"o4o]oXojo |o�o�o�o�o�o�oTYSDEBUGf����`d�pSP�_PASSfB�?,{LOG �V���`�h�  ���a
�MC:\XtYr_MPC^}������q
� ��vSA/V �a}~t�r��e�wSV|T�EM_TIME �1�� (�`v��dk�h%�T1S�VGUNS�g'�����ASK_?OPTIONf������BCCF�G ��G� @�*��`3�9A� j�U�g�����ğ��� ӟ���0�B�-�f�Q� ��u�����ү��ϯ� �,��P�;�t�_������e��ſ����
� ���@�+�d�Oψ�� ���}����������� ��B�0�R�T�fߜ� ���߮��������� >�,�b�P��t��� ��������հ�*� H�Z�l����~����� ��������2 V Dzh����� ��
@.Pv d������� �/</*/`/�x/�/ �/�/�/J/�/�/ ?&? ?J?\?n?<?�?�?�? �?�?�?�?�?�?4O"O XOFO|OjO�O�O�O�O �O�O�O__B_0_R_ T_f_�_�_�_v/�_�_ oo,o�_Po>o`o�o to�o�o�o�o�o�o :(JL^�� ���� ���6� $�Z�H�~�l������� ��Ə��� ��_8�J� h�z���
�������� ԟ
��.���R�@�v� d�������������� ��<�*�`�N�p��� ������޿̿��� �&�\�Jπ�6��Ϫ� ������j���� �F� 4�j�|ߎ�\߲ߠ��� ������
���T�B� x�f���������� ����>�,�b�P�r� t�������������
 (:L��p^�� ����� 6 $ZHjl~�� ���� //0/V/ D/z/h/�/�/�/�/�/ �/�/?
?@?��X?j? �?�?�?*?�?�?�?O��?*OFH@�$TB�CSG_GRP �2�E��  �HA 
 ?�  sO�OoO �O�O�O�O�O_�O'_�9[LBSC�ZLd�0 �hQ?HA	 wHBH9XL�̈́V>8TB   CyP�_0�[xZ�_�RD�_�]�A��_pQ�UA�QT8Q1o�Z6ff�_^ge@H@C�_�n@�^o�j	`C��o�o�o�n �_�ohVh<uO ,z�bt���{�?Y���t�	�V3.00kB	�lr2c�s	�**�"�GB9��v�a��33H@\��y 8p�B�q�  �������LAJCFG -�EdA g@��+���������5�C�@C� i�T���x�����՟�� �����/��S�>�w� b�������ѯ����� ��=�(�a�L�^��� ������߿�kB�0�� � �ʿS�>�cω�t� �Ϙ��ϼ�����+� ��O�:�s�^߃ߩ�HA 4O��O������(�� L�:�p�^������ ������� �6�$�F� H�Z���~��������� ����2 VDz ��?��`��� 
@.dRt� ��|���// </N/`/r/,/�/�/�/ �/�/�/�/??8?&? \?J?�?n?�?�?�?�? �?�?�?"OO2O4OFO |OjO�O�O�O�O�O�O �O_�6_H_Z__�_ x_�_�_�_�_�_o�_ ,o>oPobo o�oto�o �o�o�o�o�o: (^L�p��� �� ��$��H�6� l�Z�|�����Ə��� ؏���� �2�h�V� ��z���l_ڟ쟪� ��.��R�@�v�d��� ����Я������*� �N�<�r�������b� ̿���޿ �&��J� 8�n�\ϒπϢϤ϶� �������4�"�X�F� hߎ�|߲ߠ������� ��
���T�Οl�~� ��:����������� �>�,�b�t�����V� ����������(: ��p^���� ��� 6$Z H~l����� �� //D/2/T/z/ h/�/�/�/�/�/�/�� ?"?���/d?R?�?v? �?�?�?�?�?OO*O �?�?`ONO�OrO�O�O �O�O�O_�O__&_ \_J_�_n_�_�_�_�_ �_�_�_"ooFo4ojo Xozo|o�o�o�o�o�o �o0@fT� ?6?��p��� ,��P�>�t�b����� ��Ώ�������� L�^�p���<�����ʟ ���ܟ�� ��H�6� l�Z���~�����į� د���2� �V�D�f� h�z�����Կ¿��� �.��F�X�j�Ϛ� �ϾϬ��������� <�N�`�r�0ߖ߄ߺ�8������  ��� ����$�TBJOP_GR�P 2�����  ?�h�4�;��B����O0O���@�^}� � ����� ��S�	 ��BL  ��Cр� D"�S�����?�fff��:l�B ���ff@����33D   ���+�6�����h�z������9<�b�Y��?٢�������A���D��$��[�������
9��P�A��@����C�R�= ��U�A6ffhX�D/��z��͌�� ���a�9�����!@1�tz�&���{�333<T�8o���?��?L� 9 S�B�Zcu��

� >�ff�D��L^� ^�%/F8/"/0/^/ �/j/$/�/�/�/�/�/ ?�/�/>?X?B?P?~?,�?�C���1�5	V3.00���lr2c��*��0���OG �E���E�A �E��E��3�E�iNE�!h�E�فEۑ��E�I�E���E���E�r�F�F��FM(F�5�FBFaO�F�\F"f�$Bz  E�@ �E�� E�� �E�  E��@��� E��@�� �E�~@Ԇ@�~@��� F   F�� F$ Fj�` F�@ F��P F�` 9��IR9�o�<D�ED:��O
R��S�DI_0�ESTPARS�@��M��1�HRcPABLE� 1�B�,P�DNX#W |�YNWNX�NX��NW	NX
�NXNX�U�NX�NXNX�A}SRDI�_L��_�_�_�_�_�U^dOfoxk�o�o�oH�o�n~RSdoJ� (j �������	� �-�?�Q�c�u����� ����Ϗ�'�cpg�\ "�/A�_�_o�#o5oGh~R�NUM�  ��L����� �@�@~R_?CFG �񛞓���@4�IMEBF_TTiQ��J�vP3�GVER�C4�I�3��R 1�B�
 8IO�ড ��-�  ������į֯ �����0�B�T�f� x���������ҿ��� �Q�,�>�T�b�t�s��_�`�@J�
4�M�I_CHAN?� �J� ��DBGLV�I�A�J�3���ET�HERAD ?*��3��K��τ�xL�.���ROUT]�!B�!~Ԝ�o�?SNMASK(�J�>9�255.���3�����0�OOLOF/S_DIiP����ORQCTRL C�k��c_f�8U� ������������� �,�>�}�z�L�^����_QPE_DETA�I�+�PON_S�VOFF!��P_?MON ��H��2��STRTCH/K �B�eߦ��VTCOMPAT���3Ӥ���FPRO�G %B�%  ?AL_TCP5����PLAYjX��_�INST_M�� 2����US]�U�gLCK��QUICKME��!goSCRE>+�tps�0g�Y^��o_s�PR	��SR_GRP �1�B� ���.����/�3/!/W/E.�0�~/�* Q!��/�/�/�%�?? �/'??K?9?o?]?? �?�?�?�?�?�?O�?�5O#OEOkO	12?345678O�O�^RXX1��
 ��}ipnl/��@gen.htm��/�O__(_:_Pp�Panel s/etup>\}4~_`�_�_�_�_�_ m_ c_o"o4oFoXojo�_ �oo�o�o�o�o�o �o�oBTfx�� A7����,� >��b���������� Ώ��W�i��(�:�L� ^�p������ʟܟ � ����6���Z�l��~�������+��UA�LRM� G ?B�
  ͯ�� �J�=�n�a������� �����߿��4�西SEV  ���f��ECFG �����ƍ!A�� �  Bȡ
  5ϡ+���������� #�5�G�Y�k�}ߋ�r����� ��/���@�Ik?u�(% (�� �A�,�e�P� ��t���������0��+���� �����9�I_=HIST� 1���  �( c���%/�SOFTPART�/GENLINK�?current�=editpage,,1 �����0����
�(�����menu��955 ����m� 2D�148,2 _XY\����53��Z�w��*<�0f�//d,/�'�E34�����4��/�/�/�,C/��CAL���/?`"?4??/Q/��71���MV�/�?�?�?�=� !��!��?�?OO/O AO��?kO}O�O�O�O �OTO�O�O__1_C_ �Og_y_�_�_�_�_P_ b_�_	oo-o?oQo�_ uo�o�o�o�o�o^o�o );M�o�o� ������?�� %�7�I�[�m�p���� ��Ǐُ�z��!�3� E�W�i���������ß ՟������/�A�S� e�w��������ѯ� �����+�=�O�a�s� �������Ϳ߿�� �'�9�K�]�oρϓ� ������������ߠ� 5�G�Y�k�}ߏ�߳� �����������C� U�g�y���,����� ����	����?�Q�c� u�������:������� )���_q� ������� %7�[m�� �DV��/!/3/ E/�i/{/�/�/�/�/ R/�/�/??/?A?�/ �/w?�?�?�?�?�?`?��?OO+O=OOO:
��$UI_PANE�DATA 1�����A�  	�}  �frh/cgtp�/widedev.stm[O�O�O�O|�O�L)  ri�O &_A �@>_P_b_t_�_ �_�O�_�_�_�_�_o (ooLo3opo�oio�o��o�o�o�o :�� �  p # Q�8_=Oa s���o�._�� ��'�9��]�o�V� ��z���ɏ���ԏ� #�
�G�.�k�}�d���y���C���� �)�;���_������ ����˯ݯD����� 7��[�m�T���x��� ��ٿ�ҿ���3�E� ��ʟ{ύϟϱ����� (���l��/�A�S�e� w߉��ϭߔ��߸��� ���+��O�a�H�� l������R�d�� '�9�K�]�o������ ���������#�� G.k}d��� ����1U <y�������� �	//n?/��c/u/ �/�/�/�/$/�/�/�/ ?�/;?M?4?q?X?�? |?�?�?�?�?�?O%O ��[OmOO�O�O�O O�OL/�O_!_3_E_ W_i_�O�_t_�_�_�_ �_�_o�_/oAo(oeo Lo�o�o�o�o2ODO�o +=O�os� �O������j '��K�]�D���h��� ����ۏ�����5�0�Y��o�o}�j��� ��ǟٟ���)��"� �u�N�`�r������� �̯���ׯ�&�� J�1�n���g�����ȿ�ڿ�����x�c�k�$�UI_PANEL�INK 1��e�  ��  ��}12�34567890 W�i�{ύϟϱϹđr U�������)�;��� _�q߃ߕߧ߹�Q�Q��
��ݘqS�  �SOFTPART�/GEN9�?CO�NFIG=SIN�GLE&PRIM�=mainedit ��A�S�e�Q�
���M=wintpe,18�������� ���.�@�R�d���� �������������� *<N`r
�� ������&8 J\n���������� 0,�  1� E5�or
�K.- co2/s/V' �/�/�/�/�/�/�/�/ ?1??U?g?J?�?�� �ߞ?�?�=R��OO /OAOSOeOX��?�O�O �O�O�O�OxO__1_ C_U_g_���e�a�]�R �_�_�_�_�_	oo ��3oEoWoio{o�o�o .o�o�o�o�o�o ASew��*� �����+��O� a�s�������8�͏ߏ ���'���K�]�o� ��������&'ӟ�t? 	����?�"�c�u�X� ������ϯ����� )�;��4�]�_�?u_�? ����п�����O*� <�N�`�rτ�ϨϺ� �������߃_�_�_ \�n߀ߒߤ߶�=��� �����"�4�F���j� |������S����� ��0�B���f�x��� ��������a��� ,>P��t��� ��]�(: L^͟����� ���/�6/H/+/ l/~/a/�/�/�/�/G� �/k� ?��D?V?h?z? �?�?�?���?�?�?
O O.O�?ROdOvO�O�O �O�-�?��__*_ <_N_`_��_�_�_�_ �_�_m_oo&o8oJo \ono�_�o�o�o�o�o �o{o"4FXj �o������� ��0�B�T�f�x�� ������ҏ���e� ,��/P�b�E���i��� �������՟���:� L�/�p����/��?ʯ 9?� ��$�6�H�;O l�~�������ƿؿg� ��� �2�D�V��O�O �O�ϰ���������
� ��.�@�R�d�v߈�� �߾���������*� <�N�`�r���%�� ����������8�J� \�n�����!������� ����"��FXj |�����e�� �0TfI� m������/��υϿ�s-�$U�I_POSTYP�E  ��/� 	c"s/w/�_QUICKMEN  �+b/�/�!�RESTORE �1��  ��"*?<?`9m[?�?�?�?�? �?o?�?OO&O8O�? \OnO�O�O�OO?�O�O �OGO_"_4_F_X_�O |_�_�_�_�_�_y_�_ oo0oBo�OOoaoso �_�o�o�o�o�o�o ,>Pb��� ��yo���q#� L�^�p�����7���ʏ ܏� ���$�6�H�Z� l��y������؟� ��� �ßD�V�h�z� ����A�¯ԯ���
�ހ'SCRE� ?��-u1sc�%0u2E�3E�4�E�5E�6E�7E�8<E��"USER'�,�2>�T&�G�ksO���U4��5��6��7���8��� NDO_C�FG �+  �$0 � PDAT�E ����None V� S�EUFRAME � $��$�RTOL_ABRT/Ϝ�"F�ENBP�A�G�RP 1�9�!?Cz  A��ä��	!�϶�����������?�� Up���_�?MSK  s�{њ_�N,�%Y%|�%����߂"VISCA�ND_MAXq��I�[���FAILO_IMGq�^ �	 �#{���IMREG�NUMq�
���S�IZq�$0����,�ONTMOU4O�s����N��_�d � ~���¿FR:\�� �� MC:�\P�\LOG��B@�� !����������%z �MCV����UDM1(�EX1������TRAIN���^ o���)� (ޡ!=��ͧ��� ������������� "4FXj|�����PO64_7〜���&n6�I�L!I��
�V����f@�� =�	SZV����WAI��S?TAT ��	 !@�����$�/���H�2DWP  ?��P GC �"��2(9�A/��_JMPERR 1�+�
  ��2345?678901�&�� �/�/�/�/�/??8? +?\?O?�?s?�?�?�L�MLOW�����δ�_TIW��'���MPHASE � ���-@��SoHIFTM�1'��
 <�<��vOE UO{O�O�O�O�O�O�O  _�O	_/_h_?_Q_�_ u_�_�_�_�_�_o�_ oRo)o;o�o_o5E����	VSFT�1�V��M�c S�5��� �����A�  B8�`��`���psq�b�s]ЬgME> s���q�f	�&%�5A�M������1���$�TDINEND[�\؎tOp�S߬w�Y��S��y�0q����G�#��F���&��&���xRELEAqϋtV�h�q?_ACTIVԉ|�<
��A �ۗoV��
�RD� Տ�YBOX �ｬ�������2�X�190.0m.�83����'254��0A��� �(�:�����robot�d�� ?  pF�{���pcɐ�����Ꝋ�����a����ZWABC����,�  %��⚯O�5�r�Y�k� }���̿���׿�&�@�J�1�Cπ��Z9������