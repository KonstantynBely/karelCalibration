��  ë�A��*SYST�EM*��V7.7�077 2/6�/2013 A�Q  �����ABSPOS_G�RP_T   � $PARA�M  �  �ALRM_�RECOV1   $ALMO�ENB��]ON�iI M_IF1� D $ENA�BLE k LA�ST_^  d�U�K}MAX�� $LDEBU�G@  
FPC�OUPLED1� $[PP_PROCES0 � ��1��URE�Q1 � $�SOFT; T_I�D�TOTAL_�EQ� $,N�O/PS_SPI�_INDE��$�DX�SCREE�N_NAME {�SIGNj���&PK_F�I� 	$TH{KY�PANE7�  	$DUM�MY12� �3��4�GRG_S�TR1 � �$TIT�$I��1&�$�$T�$5&6&7&8&9'0''��%!'�%5'1?'1*I'1S'1]'2h"GSBN_CFG1 � 8 $CNV_JNT_* ��DATA_CM�NT�!$FLA�GSL*CHEC�K��AT_CE�LLSETUP � P� HOM�E_IO� %�:3MACROF2R�EPRO8�DRUeNCD�i2SMp5�H UTOBACK}U0 � �	�DEVIC#TI\h�$DFD��ST�0B 3$INTERVAL��DISP_UNI�T��0_DO�6E{RR�9FR_Fa��INGRES��!Y0Q_�3t4C�_WA�4�12HGX�_D�#	 d �$CARD_E�XIST�$FSSB_TYPi�� CHKBD_S�E�5AGN G�� $SLOT_�NUMZ�APRE�V��G �1_E�DIT1
 � Uh1G=H0S?@�f%$EPY�$OPc �0L�ETE_OKzBU�S�P_CRyA�$�4�FAZ0LACIwY1KR�@k �1�COMMENy@$DGV]QP� h���AL*OU�B? , $�1V$1AB0~ OL�U=R"2CAM_;1� x�f$A�TTR��@0AN�N�@�IMG_H�EIGHyAcWI7DTH�VTCYU��0F_ASPE�CyA$M@EX�P;$� Mf�C�FcD X $�GR� � S!1U`BfPNFLIC`~d
�UIREs3��AO}MqWITCH}cJX`N.0S_d�SG0� � 
$WARNM'@f��@� sLI? �aNST� �CORN��1FL{TR�eTRAT@0�T�`  $ACC�1"p '|�'r�ORIkP�C�kRT�q0_SF� �!CHuGI1 [ �Tz`u3IPpTYPVD�@*2 �P�`�� 1zB*HD�SJ�* ��q2�v3�v4��v5�v6�v7�v8��v9�vqO�$ <� so�o�h�s1��PO_MOR._ t 0Ev�NG�8`TBA � 5c���A�����]@B����ϋP�0XЅ*��h�`
P@�@�2� �,p�J,pC_Rrrqo@+�J/rL/�J�JVq@�Cj�`�m�g��ustP_}0sOF� 2  @� �RO_���WaIT<8C��NOM_�0�1�ەq3� ��cD !�;����hP���mCEXpG�0� F�<p%r
$TFx�J6F�D3ԐTO�3&@yU=0�� �YH�24�T1��E�� �e��f��f�>�0CPDBG;a� mk@$�PPU�3�f):��A��AX 1�dUN�$AI�3BUFuF��⠎�! |�`��`P�I��Pr�M�q�M~�䠁�Fr�SIMQS��G��Q�E�����MC{�5 �$}1JB�`S��}1DEC��������ܴz� ě0CH�NS_EMP�r#$Gg�=Ǎ@_��q3�
p1_FP󔞡TCh�@`�b��q0�c}�y�G�� V�AԂ�!!���JR!0ԂSEGGFRA.pv 7aR��T_LIN�C��PCVF������Y ���Q��)B����( '���f�e �S���Q��.0�p�B�8�A����SIZC����z�T��g������QRSINF3��p�� ��?�������؉����Lot��G�*�CRC�eFCCC�`+���T� h��mh�SbA��h�*��f��:�D�d�c��C��PTA����w@��L����EV���jF��_��F��N&�G�� �X������1i��! ��,��h#RGNP��0qF���R�}�D���2}�LEW N��Hc6���C�K���}RcDx :�@L��ou2���A6N`�Co�$LGp��B@�1aP��s@�dWaA?@����~0R���dM�E%`��d�_RAs3dAZC���z��OkqFC�RH`X`F�`��}��,�ADI ;� 6b� ���` �p�`5cn�S�@1�L7a�AMP���PY8C�U�MwpU��iQU� $�P��C�C�G1������DBP�XWO����p�$SK��2� D�BT TRL�1 ���Q0Ti� �P�D�J�4LAY_CA�L�1R !'PL	3&@�0ED�Q5'�Q�5'̡PP���1!��W�PR� 
p�1 0�1" �P�A$�q$�� �L�)#�/�#mpR�0$�/�$C�!%�/��$ENEqr�&��/�#d REp�"'�H �O)@7"$LF3#$�#xBП W;���FO[ _D0m�RO(@���u���j���3RIGGE�R�6PA%S���E�TURN�2RcMR-_��TU�`?�u0�EWM����GN�P��zBLA��E��/$$P#�CP� "��&@�Qk�C5D�mpD�A#�p4\1i�FGO_AWAY�2�MO��fQg�C�S_(<�QIS ����c�C���A����B�t�Cn�ȫA"�FW���DNT	V@��BVkQ�����S˳W�sU�J&�U�� ���SAFE�ZV_�SV6bEXCLUtl�����ONLA�b�SY��Q�tOTBa���HI_V/M�P�PLY_�a��VRFY_#�q�Bd��_ )0���_�+�Ip ���ASG3� *�b݀�0  AA��a*����0���Vi.b%fANNU�N� rLdIDp�U�2~S@�`mijaprj�f�pOGI�"+��$FOb�׀�OT@w1 $DUMMY���d[!��d١�& �E, 7` 8�HExs���b�SB$�SUFFI�@ ��@�a5�g6�a!�DwMSW�E- 8���KEYI����TM`Z1^ӌq�1�vIN��⎀�. D޵�HOST? ! �r���t[ �t٠�tYp��pEM>���$��S�BL��UL��/ A�|3����T50~�!0 � $9��ESAMP�ԕF��������I�0��$SUBe�Q�� ��C�:��G�SAV ��r���G�C� ˇ�P�nfP$80E��YwN_B�1 0��DIad�@O���}�$]�R_I��� �ENC2_S�T � 2
ԇ J����L�q~S�`;����!3��M�I��1:�p�4  L�3�M��0��0K�4'a��AV�ER�q��}�M�DSP�v��PC�U����\ì�VALU�ŗHE� ��M�I�P@���OPP7  ��THS ���6�SH�F�F􁳠dL��0�T��SC�Q�d�:�ETo�5zrF?ULL_DUY�da��0��O�w�h�OT����0NOAUT5O�!6�p$�\֤��cl�
�C` ��C���`!�L��� 7H *��L���n�b���$ �0P�˴��ֲ��[!��@�a��Yq��dq��7���8��9��0����1���1��1��1Ⱥ1�պ1�1�1��2R
�2����2��2��U2Ⱥ2պ2�2�U2��3
�3��3�����3��3Ⱥ3պ3*�3�3��4
��Qv��SE�"8 <��~��`�;I����׌/��QFE�0�0� 9� ,��Q? �z@^ ?�А���ER@#�,���A��� :�`$T�P�$VARI�� �s��0P2�P; �pq�TD��S|��1`3���e�BAC�< T�pr���)��bP�P o�IF�I)�P ���U���P�� ��0��� =t ;'�Ԡ��P'�ST(&�� HR&�Pr0E����	%�C��	���_Cr�N�r��B���p�h�FORCE�UP%bn�FLUS
�`HN �E�h�R/D_CMK@E(����IN_��&vPg�REMM�F~Q���M �� 3
K	N0�EFF��N@sIN�A��OVMl	�OVAl	TROV̙��DT��mDTMX���m{@�
���? �*[ ��CL���_:p']@$�-	_�
�;_T��X
�J�@AQD� ��}���}!V1� RQ~��LIMIT_�ad椀�M��CLmd�}�RIV	�a��E�AR��IO*PC�C�����B�Bg�CM�@��R �GC3LF�G!DYM(/l�aR#5TWDG��h| s% �SS& �s> P�a�!r1��EwP_�!�(�!1���E�3�!3�+5�&��GRA���?w�4�kPW��ONT��EBUG)S&2*�P�{@a�_E @ ��p�R �TERuMB5AK9ORI�G0BK5�`�SM_��Pr�G0CK6U0A��9DK6 �UP>B�E� -zAa��@.PY3.@A$S�EG�:f ELEUU�SE�@NFI,���2�1ޠp4�4B$sUF6P�$��FQ4@�wAG0T�Q�&�HSNST P�ATm�piBPTH	J�AߠE�p��2�P@؀	E)�؁��1R�@<�InaSHFT_��1|oA�H_SHOR �ܣ�6 �0$�7�@Dq�'�OVR#�na�@�I�@�U�b �QAGYLO=�z��I'"��oAj�!�j�ERV ��:Qh��J��OG @�B�0����U>���R!P"�ASYM.�"��1#WJG�уES�A�YvR�U�T @���E)�ᥳEP!�WP!�W�OR @MB��GR�SMT�F�GR��3laPA.@��`|�q�uG � ����TOC�1�`P<�@ �$OP���P�pՓá ��O�񖌀RE�`RC�AOX�pтpBe�`RmE� u�h�A��e$PW�R�IM�ekRR_p�c4��qB H2�H���p_ADDR~��H_LENGqBPyqnq�q�R��S�I H��S���q0���u>Ӵu���u��SEȸ'�LrS��J� $��`��_OF�F��rPRM� �Z�HTTPu_�H�K (^p�OBJ?"ip��$���LE`C!�ȠL� � �׬�AB%_~TS�s�S{`��6*�LVN�KR��e�HIT��BG��LO�qt�fN�͂���`���`SS{ ��HQW��A�M�p`�INCPU�"VISIO�����+��t�,��t,��� �IO�LN��N̠�C^��$SLQb��oPUT_�$�`�{�P �W���F�_AS�"O��$AL��I����A��U�0��@Af��`q�<PH�Y���Ó�ў�UO��#P `�����@�ڔ� �2�pP���`(�L��Y�B���UeJ�Q�z�NEW�JOG-G��DIS�x�[�K-�f�#R �
�WAV�ǢCTR<�CǢFLAG�"[�;LG�dS ����Y�3LG_SIZ�o���������FD)�I�4�E�*�� D0���c$���𖶀����K���D0��� SCH_��߅p�2���N��F�T���E �"~�������U
�
�r{`L�	�DAU/ŃEA�-��dE�;�G�H�b�OGBO}O��Uh Aɒ���IT��y�[0ŖR;EC��SCR�𙃖ʑDIēS.@��RGO���˒����d��$����SU���W�Ĳ��Ľ�JGM$�MN�CH,�FNKEuY%�KM�PRGK��UFY�PY�FWDvY�HL��STPY��VY�@Y؀�Y�RS"��H1`uۺ�CT�� �R��� �$�U	�m�@��
R�ݠғ`�G=ن�@POd�ڻŦ�M��FOCUd�RG�EX��TUIK�I{�����	������I�M��@A�S�`��p�@������ANA����2�VAILl�C�L!�UDCS_H!I+4`�s_�Oe�
!"h�S���|�S����IGN4��F�J��9T�be�_BUj � �V !PT�$�*��rv�ϤS1��A
VrW !Pi�'��T�0�1?2?3?�!��`� X � �i�=a�5���Ņ�IID� tbP5R�bOh X��\A�ST	�RF��Y�0�@�  W$E�C�y�����_�� Y L �؟0��@���`q�Ftǀ�FwҬ�_ Z �p����b���>0C��[ ��p CLDP	��UTRQLI{��T����FLG�� 1�bO�D�����LD���ORG����� �hW>(�siT�r� 4\ �#0��վ�%Sy`T�70#0' ��$�!�#RCLMC��$B/T/�)Q��!=1I��p_d] d�R}Q73$DSTB�pƢ   6��-8AX��R /8I<EXC#ES�bd�2Mp�1�^�12�Tt6��0_�p"6_A:&��;�G?Y80K�d` \��GROU��t$�MB �LI9�CREQUIRDB�aL=O#KDEBUr� 1LYM��agbʑ`@h�C�" 1ND���`c`b���̨�CDC���IN'��C��Z`���H��N�"�a#�� �EPST�� �c\rLOC�R!ITp��P�Ap��1 1ODAQ��d� X�ON�cF �R�fV�	X��b�U����w �FX0I�GG�� e ��y X�a��X�XR�Q%��Y	��X	�x�V�0ғDATAB$`E�a��a�N���f t $MD
EaI:�)Sf��^d�![gH5P�@]ez��a_cANSW�a^d�a��
^eD�)ARz�� Xp�g �0CU4�V��`�=URR2{�h� D2�`A��A�! d$CALI&0ү�GS�w2K�RI�Nb�t<�NTEg�(i�bCu��=RBqg�_N�qjPukr����$ht�2kuyDIVF�&DHi0jp+�l �$Vp�C�$M�$Z0R<!T 0R����b�emH ?�$BELT˪Z_ACCEL���;�"�IRCO�݁m���T���$PSi0�L ڰW���Cp8��T�9�PAT!H���.���3]��Pl1_<�r��Ł�"S �Cr��_MG���$DD�9���$FW�`7`���.����DE�PPAB�Ne�ROTSPE!EՂ@L� JN�@�(0� $US�E_p�P&�ܦS�Y>��p�! �QYNr0A����OFFuan��MOU߁NGJ��܀OL~�ٔINC �d2Q��-2��� -2ENCSpa2U�X�+4R�IN�I]�0B����"n�VE��s>^�23_UPօp�/LOWL��[�` '���D>�2@Ep�]'��2C[pW�MOS���4MO��0�'PERCH  ��OV����蓼��� ���$�8S+�� 2@�������V�0^�O�L`�P��7O�U�UP"�8������TRK��AYLOA�J��1���]�͵³3P� �RcTI�1	�� MO� O�-2�28 �`4�w�ٳ��?�pDUM�2��S_BCKLSH_C]�P�ϐΦ ����bn�"�y�Ñ���CLAL V��!8��� ��CHK �SՐRTY����C��
*!6a_�ä_U�M����C���SC�L�W�LMT_J'1_L< 0-օa:�E4�U�G�D�J�P�J�SPCd�ȑZ���&3�PC �3�H_A@d���C� cXT��.�CN_rN���".�S��%�V���@:����]�9���C' �SH�r�*�*! 9�9� p��^���9���3PA���_P��_�"�Ŷ�!ճ�����JG����~�OG|��,�TORQU��ON��޹*�B٢-�L*�L�_Wž�_�s�j��sj��sj�Ir�IJ��I�sFKP]�J�!X��c!�VC�0'42��1��{0��82���JRK��+� D�BL_SM���"Mζ@_DL�q�"GR�Vq�j�sj�sKH�_��I���
COS��LN- ��� ��p�	�p�	���ĺ�FZ� ٦KMY��D�TH�eT�HET0��NK2a3�s��s� CB�CB�sC&1n2���0��s��SB�s�N�GTS�1W�C.� 2Q�����$�'3$DU���8A!r �2P&�1Qb8V'$NE�4�PI� ��H�"%�v$�p�A��%�'���LPH�5�"h��"S��3� 33�"+3:2�pEV�(V�(�p�,V�*UV;V;V";V0;V>;VL9H�(�&�2P�-n�H;H;H";UH0;H>;HL9O�,�O�(O}I�.O�*O�;O;O";O0;O
>;O2F�"�Y��T�'SPBALA�NCE_T@SLE6�H_�SPHq��hR�hR3PFUL�ClX�R{W�R3Uz1=i
�UTO_�����T1T2�Y�2N ���`��Tq���Ps (d���T�O�p!�>L�INSEG����REVf��Q�DI�F��zy1j_g�r1k��OBUa��t$y�MI`���SLCHgWAR>��AB��~u$MECH��Tˑ�a��AX˱P�y��f�'�r�Pl 
p�bI��:�ROB㠣CRW�-u�Ҕ�pM�SK_KP�tn P+ �P_��R��r_tn���18�c�a�_p�`�y�_p�aIN:a��MTCOM_C|���po  ݀�g`4�$NORE�S��r��`�rp �8U�GRJ��eSD�� ABג$XY�Z_DA�!F�r�D�EBU:a�q���pqu _P$��COD��G 1����`���$BUFIND�Xa�Hp"�MOR^Rsr $�qU&� ��u��ӑy�^��b�Gi�s � $SIMUL��8��x>���F�OBJEjP>��ADJUSψOAY_I��8�D����s�Ԑ_FIב=s�TZ��c�����`b�"�(�b`p0G�DN��FRIW�d�Tg�RO%�A�Eb�}П�OPWO> Vpt�0>�SYSBU<0[�$SOP��I�����U��b`PRUYN�rڕPArpDٖ��b��1�_OUT�Α�a�t$�IMKAG��\pv PDa3IM��1�IN[ �~0�RGOVRDY�˒���P�/�a�� �L_�PB�}����R)B�� ��MkᜪSEDb��` �N�@�M��~�Hp\�SL�jPVpu x $�OVSLfSDI��DEX���q����H�o��Vb��N��A��'��,�'�D�M�~Ҥ_SETK�Vpv @U�^��e�p�RI��j�
q�_�}�����Hpdà>*� w H\q�`���ATUS<�$�TRCx T�X�ѳBSTMڷıI��P��4}Ѱ���Vpx DB\pE���β�0Ehb�ϱ�����ϱEXE�հ����)�=��f�y�m�]p԰UP�L�9$�`6�XNN����x������ �PG�u7zWUBñ�e���ñ��JMPWAeI[�P���LO7���pFA`��$RCVFAIL_Cwq�p��R9��p�c��(��}�"�-�AR_PL��DBTB��,��pgBWD ��pUM*��"�IG�7��Qc�T#NLW�"�}�Ry�iӂ��E�����Hp��D�EFSP` {# L\p�`��_��Ճ��UNI����Ѐ��RD��Rb _LA`PJͱ��P�pUq|-��#��q�O��XPc�NN�PKET�
��Pq�Uq} h�ARSIZE5p��=���u�S̀OR��F�ORMAT�Pg�C�Oנq�<bEM�d�����UX��,�5p��PLIb�Uq~ � $�pP_SW�I�`��/ G�b�ALO_ o���A�r�B���C�rD���$EL���C_�lі� � � 1���r��J30 �r^��TIA4Z�5Z�6�rMOM��f���s���pB��AD`f��s����PU�NR����s���������Rt�� A$PI�&E�kqE�p- ~-�-�WC�0$��&�9q�gE���eSPEEDL@G �����Ծ����)� 9����)��	)���SAMWPx�0�1��MOVD�H$_S` Y%nk%_��1�t�2�t����c�v��8�H�PxIN��� ������(�+(+GAMM<Vu!�$GETE�U�ٓ�D5�
�PLIB�Rv���I�$HIBu�_L�ݰpB�&E�b�(A�.� �&LW�- �&�,�)	6�&1��f�`�j��� $PGDCK���ٓ_�����E���b7���a4��a9�� W$I��R�`D�c0�b~�Ե`LE�qkq��81��0�,���`Vp�P/aUR_SCR��A�r���S_SAVE_�D��8Ex�NO5�C ��y�6�8@{$E�.{I ��G	{I�@�J�KP�q ��H� ���x"Ma o���s����d� �6W2U�Cqy�ѡ��M� �k�F�� aE��3�W<�@[�jQ!Wg@5r�U�R�R��ȥSc2jQM"��[CL��W��M)ATr� �� $PY����3$W`�fNG�O� `�b�b�b#�HЈ��a� ���c��X�O���Z�e��ހ�Rt� p䠰p�3 +zO�O�O�O�O�a5�_�r� |�E�8@ ��>vs�>v��8@_�kwVvy�Eހu%�!sB��\�P�"tP����PM&�QU5 �� 8*�QCOUܒ1 �QTH#pHO�L<�QHYS��ESe�qUE�p.BZ�]O��  q�P��̕%��UNְ�Q ���OE��p� P�2�3��AÔ�ROQG�����Q2(�O}��2������INFO�q� #�e����R�Ⱦ�OI��� (�0SLEQ�с��рi�C�{�D��L��D`� OK0r��!�E� NU!��AUyTTA�COPYqPu�?��`@ML�NI��M�X�Cᐛ� Y�R�GADJ�q�i�X�Q��$ഖ�`��W��P���0��������EX8�YC0b$�ѪObp�q���$�7_NA9!��������`��� �s Q���PORӸA�B�SRV0�)la�Y�DI��T_�� {�������������U5��6��7��8y�Ҿ�S8BL��m�MCS_F�p��PL9A8An�ȰR��9��Ѽ���$iB����d� �,�0FL-`L�C@Y�N�[�M��C?��GPWRc��L��!�ODELA��8Y5��AD�a��QSwKIP� �Q�Z4�OR`NT�Q ��P_4��ַ@lb Yp������ ����Ƞ��ՠ���������9�1�J2Rܻ L�� 4*�EXs TQ%����(Q�����p�����p���RD�Cf� �`��X9�R�p�����r��~A$RGEAR_� sIOT�2FLG��vi��M%PC��B�U�M_����J2TH�2N'�� 1������G8 T00 I�����MlѺ`I�\8�qREFr1�q� l�h��ENA9B{�(cTPE�0� 1���i�m���^QB#���:��"������2�ҙ����������
&�3�Қ7�I�[�m�(��&�4�қ�����������&�5�Ҝ�1�C�U�g�y���&�6�ҝ����������
&�7�Ҟ+=Oa(s�&�8�ҟ������&�SMS�K�q�|��a��E�?A��MOTEF����a@��(Q�IOQ5�Ic(P�Pά�POW�0L�� �pZ����#p%�L���U�"$DSB_SIGN�1)Q%���yCl��S232���b�iDEVIC�EUS�,R'RPA�RIT��D!OPB�IT`QY�OWCONTR;�(Q��O�'RCU� MDSUX/TASKT3N�p[0ހ$TATU`P�V"�0L����p_�,PC9�$FRE?EFROMSp���%�GET�0�UPeD(�A�2��SP� �J��� !)$USA^���6���ERIO�P@bp�RY�5:"_>@ �P8}1�!�6WRKI[�D���6��aFRI�ENDmQ�P$U�Fw���0TOOL�FMY�t$LENGTH_VTl��FIR�`-C�RSE<N ;IUFINR]���RGI�1ӐA'ITI��4GXӱCI6�FG2�7G1����3�B�GPR� A��O_~ +0!�1RE`Ѐ�E3�e�TC��8�Q�AV �G8��"
J���u1~! ��J �8�%��%m��5�0>G4�X _0)�L|�T�3H6��8��(�%r4E3GU�W�P�W	�R�TD����T��`а��Q�Tm�$V 2����1���9�1�8�02�;2/k3�;3�:iva�9=i�a`a�^S�jR$V��
SBV�EV'�SBQ�B
K�����&c�p���F�"{�@�2q�PS�E��$.rRC���o$AŠFwPR��Gv]U�cS'�� 7�sA6I�� 0�@DqV`��p�d`���PE0�@��=�
B5S!/� ��aRg�����R�6�N AX�!$�A�0L(A���r/THIC�1Y���h�t1TFEI��q�u�IF_CH�3�qI0�G�a�pG1bxf�з�m���S@��_J�F��PR�ֱ�S���Ԁ�d �$�SР�Z�GROU��̃TOT�t̃D;SP�JOG���#&��_P��"O������j��&KEP(�I�R����@M�R@�A	P�Qn�E^�`�!�[��SYS6��"[�PGu�BRK�B �.��pIq�p��M���΂��`AD�!̃9�BS�OC׆�NӕDU�MMY14�p@S}V�PDE_OP�#�SFSPD_OVR=���C����OR�CNm0�F�.����OV��SFR��pU���Fn��!#�p�C��A�"LCH�����РOV�s0��Wb�@M��ĥ:�RO�#�ߑ�_�p�� @�@�u@VER�ps0O�FSu@CV? �2WD6���2�ߑj2Y����TR�!���E_�FDOY�MB_CiM�D�B�BL�b>�f��attV"Q�240�/p��N�Gg�z�AM�x�Z�0���¿_M�~��"7����8$C�A�7�D����HcBK81��IO�5q���QPPAʀ=�"�M�5�͵���DVC_DBxC~� � 3"�Т�!��1�����3����pН�*���U�3��CAB ��2VӆPѣIP��c��O��UX�SUB'CPU�r	�S�P  P���90^SQ׹c��."~��$HW_C�А���S��cA�A�pl_$UNIT��l��ATTRI"���	��CYCL��NEC�A��J�FLTR_2_FI_�G(��9&��1LP�?�>�_S�CT�CF_��F_��6��FS8!����CHA�1�wᇲ�"v�RSD�4"�����q�_T��PROX��>�� EMy_ܠr��8d��a d���a��DIb0!�RAOILAC��9RM��CLOÐ C��Q*q���3q���PR��S�Q�pU�Cr�s 	��FUNC��@rRIN'PѸ0��u��!3RA��B ����8F�Ğ�WAR~���#BLQ����A��������DA����	����LD)0��Q1�q2��*q1TI2rQ�ǁ�p$xPRIA�1�"AFB�P�!�|ߠ�<`�R���MsOI��A�DF_&@؅�51��LM��FAށ@HRDY�4ORG6 H���A�0 �MULSE&@"�Q��a �G�	���m��$d$�1$1 ���0��߮� xm�EG0�̃�`ARހ���09�2o��z�A�XE�ROB�Wd�A��_�œSY������S�WRI�@s1��STR��� ��(�E�� !	%1��AB( �/&�a�ӰOT0v^�	$ߠARY�s�f"���S@	�FI���*�$LINK(���!�a_%#��%{q�"XYZp82�*�q�#OFF��R�"�"�(j Bဂj�4С��n�3FI��%7�q���j����_J���%��#�QO�P_>$H+5�3�PT�B\1�2C��i�D�U�&62�TURN��2r�5t!}��p��|7FL�`���m�0��%+*7�	� 1��. K�M�&8�2�Q�2rQ�#�ORQ ��G��-(�+p��z��� 3q�E"��T�GOV�@-A��M*�y�4 �E:�E@�FW�J� �G���D��o�*� � �A7�P��y��E�A�G`ZU:ZU�CG�ER�
��	6�E���B�TAFQ��)4����r'�AXУa2.q �c�W�c�W�c�W�p�Z �0�Z�0�Z%@�ZK@�Z ��Z
!�V� �Y� 
i � i� *i� :i� Ji � Zi� ji� zi�a�ioDEBU{�$v� u��;q��"F7O�n�CAB��6��CV�z� 
fr����u kњw�!�w�!�w�1�w �1�w%A�wKA�w��p\0��"3LAB"2�|EwЄ�҂�3 �� EERVEN�� � $q�_�NAǁ!_�PO�����` f�SN�_�MRA��� d � T���ERR�����~ TYi��RI��V"0�S��TOQ��T)PL��T�Ѕ�L�G�CJ � �p�PTl X���_VA1�b�Q���#�2�!2+�����/@��p���5�$W��V���VN�[�$�@�� ��S���Q�	EHE�LL_CFGN�� 5%�B_BAS��SRvp0�K� �S��JϐU1a�%Α2�3�U4�5�6�7�8�RO���� f� NL:�3ABn��АACKwv��)��o�u0iႩ_P�U2�COq��OU��P��ӕ������TP�_KAR��0��REm�� P8����QUE٩����@���CSTOPI_ALzs��� �p��TĠ�� SEM[�dw�k�Mw�y�TY��3SO`��DI����p��=�װ_TMKӟMANRQζ� E���$KEYSWITCH��Ѱ���HE��BEAT4���EpLE����
&�U��Fd�����S_O_HOM� O��7REF�@PRi��R(� ��C@�O0�p �ECO���� _I�OCM�4M�k�p����'�O� D�!$ۧH�U��;�M7�<�@�3FORCߣ�����OMq � Q@Etxk�U#PoQ1B�O�o3B�4x�_�SNPX_A�S��� 0ݐAD�D��(�$SIZ>ߡ$VAR��TIPr�q�G�A(ҷ��
�˨r�t�n�SV�XC����F'RIF�R��S%�7�x���NFѲEАO�� x�PSIڂTqEC*�%CSGL=�	T�"�0&�V�D���>�STMT
�o�P�\�BW�@?�SHsOWw��P�SV� �K�� ���A00�0�Q��K���O���_���i���5��6���7��8��9��A ����6������20��F��
 ����U �� ��� ����0�� �J@T��:�1G�1T�1a�U1n�1{�1��2��U2��2��2��2��U2�2�2 �2-�U2:�2G�2T�2a�U2n�2{�2��3��U3��3��3��3��U3�3�3 �3-�U3:�3G�3T�3a�U3n�3{�3��45U4��4��4��4��U4�4�4 �4-�U4:�4G�4T�4a�U4n�4{�4��55U5��5��5��5��U5�5�5 �5-�U5:�5G�5T�5a�U5n�5{�5��65U6��6��6��6��U6�6�6 �6-�U6:�6G�6T�6a�U6n�6{�6��75U7��7��7��7��U7�7�7 �7-�U7:�7G�7T�7a�U7n�7{�7��M��VP$�UPD��  �P���x��YSLO��� � ��հ�����Q�TAS�sTƠ��AL1U}U����CU��W=FdQID_Lѳ�U�HI�ZI�$FI�LE_Σ�T�$�u�_VSA��� h���+`E_BLCK�(�8bg�AhD_CPUQi��Qi���Sodx_R1�ɢR ��g
PW,�d� �aLA�S���c�a�dRUN5��a�d�a�d���5��a�d�a�d ��T�pACC����X -$&qLE�N~�3t��&p����I�ѱ
�LOW_AXMI(�F1&q�T2mwAM��ɢ����I��8��Q�yTOR.�&p�{DW��s�LAC�E���&p�����_�MAuйv�u�w�qT#CV�|��wTڱ� ;�1�<ѷt��_��s��IJ����M��ӠJ�����u���u2q2���������s�pJK�цVK~�か��3fՃJ0���JJ�;JJ��AAL��(���4�5Xr;��N1B�N��	��tL�p_k�����"p���� `5`GRO�U�PY�ӲB$�NF�LIC�ө�REQ�UIREv�EBU`V�"q���кp2����#pɖ!qxг�� �\��APPRՐC����p
!�EN�CsLOz�,�S_M �ȋ�A��u
!q��� 䣠MC�r;�XrN|�_MGц�C���,`��N��p��BRK���NOL������Rϰ_LI��է����	JޠѤP��p��p@���p;��pD��p6��K��8������� ҒMr:qxl�Gqz�PATHv��������Rx������6�pCNR�CA��էl���IN%rUC�p�wQ�Cd�UM�Yop�����QE:p�Gp������PAYLO�AͧJ2LHPR_ANqQ�L�`[�W��K�g���R_F2LgSHRё�LO\��䱕����ACRL_�����޷C�Xr9H�P"�$H��үFLEX� qJ>%u� :2Dv �p4�K�GYq�pPbt|F1Kљխ׃� ������E�� ��/�A�S�e�w��� ��y���ф���蘏��H��J�ÊT���X�� ��υ ��څ��[�� ��
�� �)��;�D��V�h�z�Y�J��� � �������QIPcAT��ё��EL4�S �ؘJ���ߐ;JE��CTRޱ���TN��F�ɗHA_ND_VBp��ܹP`�� $&�F2���K��ШRSW���Y�j��� $$	M��}�R��E��Uw�H��sA�PH�����Q���A���P��A���Aɫ���j`��D*��DɫP��G�`1)CST��9!��9!N̨DY�`���|�Y� 鰋�KыǦ�J�ч�s�U�ХP��&�/��8�A�J�S�=��� ; �t�.R66N�/QOASYM����Ґ¹���Խ��ٿ_SH�����筈4��+�=�O�JV��h�p'CI����_VI��dHN�u@V_UN!I�ÉD���J҅�B �%�B�̦D�ųD�F�̀���������*Uc����<�H�`���XQEN� v�D�IɠS�OwT�+9�XQ��� ��I�1A��äQ�`Bc��S`�  p�a.a� �� ME�����R'R�1TkPPT@�0) ���Qz�~����0�Xa	iT@�� $DUMMY}1��$PS_�ЛRF��  ��Pf6�aLA��YP�jb��S$GLB_T >mU�e�PpQ p����Q� X	�ɗ`�SuT��ߐSBR���M21_V��8$_SV_ER��OÐL�c�cCL�`�bA5��O�RTPT O�P �� D �`OB���LO˰&uq9cp�`r�0�SYSq�ADR�TP�PTC}Hb � ,&����W_NA����tz�9SR���l =��M �u`�ys�u~�s� �s���������� �0�)�T�"�5�~� ��B����s�?�?�?D>Y�XSCRE)�p5�ȐST[�s#}�P!��tX�r u_� Aq� T	� �`ob��a`�l��ҤԊ�g�c�O� ISb�c��TX�UE�TG� �ñjp^`Sq��RSM_iqmUU?NEXCEPlV֑XPS_�a����޳�p���޳R�COU�ҒS� 1�d�U�E�tҘR�b9�PR�OGM� FL�7$CU�`PO?Q��ִ�I_�PH�� �� 8џ�_HE�P�����PRY ?��`Ab_�?dGbOUS�� �� @�`v$BU�TT�RV`��CO�LUM��U3�SE�RVx��PANEԋ q��P@GE�U�<�F���q)$�HELPB�l2ETER��)_��m�A m���l���l�0l�0�l�0Q�INf��S�@N0�� ǧ1�����ޠ �)�L�Nkr� ��`T�_�B���$H�b T�EX�*��ja>�RELV��DIP>�P�j"�M�M3�?,iŠ0ðN�jae���U�SRVIEWq�S <�`�PU�P�NFI� ��FOC�UP��PRIa0�m@`(Q��TRIP>zqm�UNP�T�� f0��mUWA�RNlU��SRTO�L�u���3�O�3ORN3�RAU��6�TK�vw�VI�͑�U� $�V�PATH��V�CwACH�LOG����LIM�B���xv���HOST�r�!�R��R<�OB�OT�s��IM�� gdSX`} 2����a����a��VCPU_A�VAILeb��EX
��!W1N��=�>f10?e1?e1 n�S���; $BACKLAS��u�n���p��  fPC�3��@$TOOL�t$�n�_JMPd� yݽ��U$SS�C<6��SHIF ��S�P`V��tĐG�yR+�P�OSUR�=W�PRADI��P���_cb���|a�Q�zr|�LU�A$O�UTPUT_BMc�J�IM���2��=@�zr��TIL��SC	OL��C����ҭ� Һ�����������o�od5�?��Ȧ2$ƢN�VVp�U���vy�DJU2��� �WAITU����n����%��NE>u�YB�O� �� c$UPvtfaSB�	wTPE/�NEC�р� �ؐ�`0�R�6�(�Q��� ش�SBL�TM[��q��9p����.p�OP��M�ASf�_DO�r
dATZpD�J����|Zp�DELAYng�JOذ��q�3� ���v0��vx��,d9pY_���	�7"\���|�rP? O��ZABC�u� П�c"�ӛ�
N��$�$C��������!X`N�� � VI�RT���/� ABS�f�u�1 �%�� < �!�/�/??0? B?T?f?x?�?�?�?�? �?�?�?OO,O>OPO bOtO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_�_�_�_�_�_ o o$o6oHoZolo~o�o �o�o�o�o�o�o{� >��AXLMT�s���#  �tIqN&8qtPREO���+vupXuLAR�MRECOV ��)XrzujF }�%�!d�������7�I�[�m�~�, �
�/��vNG5� ��+	 =#��
ڏ�� PPLIMC5�?�%upՁ�Handl�ingTool �-� 
V7.7�0P/36 ���
]�_SW2�D�Fy0j�W� 43Y��J�9�K�7DA7�?����
&�X�e�	-�None���J����� �T7o�	�rP_��Viu�6s��UT�Oz"�,tTy.�HGAPON� %��!.��U��D 1�y� t�x�����y.��K�Q 1�{  THp������	��p�uq��"�"� �!��H�եw��HTTHKY��"ٯ���� u�����󿽿Ͽ��� ��)�;�M�_�qσ� ���Ϲ��������� %�7�I�[�m�ߑ��� �����������!�3� E�W�i�{������� ��������/�A�S� e�w������������� ��+=Oas ������� '9K]o�� ������/#/ 5/G/Y/k/}/�/�/�/ �/�/�/�/??1?C? U?g?y?�?�?�?�?�? �?�?	OO-O?OQOcO uO�O�O�O�O�O�O�Ƹ�TOĀ��DO?_CLEAND����{SNM  ɋ����_�_�_�_o��_DSPDRYR�_&��HI!��]@�_}o �o�o�o�o�o�o�o�1CU��MAX@ �bTQNQS�sqXbT�B�o�B���PLUG�Gb�cWo��PRC*4`B�P]klo^��rO�r=o��SEGF;�K�+�6��_�_�}�������ŏ�0�LAPZom�/��+�=� O�a�s���������͟�ߟ�6�TOTAL��v�y6�USENU
Z�g� HXL�NR���RG_STRIN�G 13�
��M,�S�
~��_ITEM1��  n󝬯��Я� ����*�<�N�`�r� ��������̿޿���I/O SI�GNAL��T�ryout Mo{de��InpB��Simulate�d��OutT��OVERRW` �= 100��I?n cyclHŕ��Prog Ab�or^Õ�>�St�atus��	Heartbeat���MH Faul<����Aler��� ��'�9�K�]�o߁��ߥ� ^S��^Q ��������,�>�P� b�t��������������(�:���WOR9���r���L����� ��������*< N`r�������PO���� ���9K]o�� ������/#/�5/G/Y/k/}/�/DEV� -�/�/�/ ??)?;?M?_?q?�? �?�?�?�?�?�?OO|%O7OPALT�� ^A��8O�O�O�O�O�O �O�O__(_:_L_^_�p_�_�_�_�_�_LOGRIxp��avO�_*o <oNo`oro�o�o�o�o �o�o�o&8J\n�_*�R�ݦqo ������(�:� L�^�p���������ʏ�܏� ���PREGbNK��$�r����� ����̟ޟ���&� 8�J�\�n���������~��$ARG_r��D ?	������� � 	$�	[�]���.���SBN_CONF�IG ��L��K�F�CII_S�AVE  ��k�b��TCELL�SETUP ���%  OME_�IO��%MO�V_H��¿ȿRE�P�|��UTOB�ACK��V�FRA:\8�� �8���'`��8�c�,�INI�a@8�^�,�MESSAGz�����|���ODE_D���}�C���O� ��,�P�AUS!��� ((O��J�\� F�|�jߠߎ��߲��� ������B�0�f�t��%�*TSK  �5ݒϕ�/�UPDT�����d����XS�CRDCFG 1v��� �������&�8�J�\�n� ��\�n���������� "��F��j|�����/e�2�G�ROUN����U�P_NAܰ��	�2��_ED��1�
��
 �%-BCKEDT-�0�}��p��ѲQ-2�p8�/�/�8���g2���E/��/��/~/��ED3n/&/�/J/�\.�/"?�/�/ED4 ?�/?�/\.[?�?5?G?ED5�?n?#O�?�\.�?jO�?�?ED6 ZOO�O6O\.�O_}O�OED7�O�Ok_�O�\.G_�_!_3_ED8�_�o�]-�_Vo�_�_ED9Fo�_�o�"o]-�o�oio{oCRoY_Vh�]1��{� LNO_D�ELGE_U�NUSE	LA�L_OUT �V��WD_AB�OR���~�5�IT_R_RTN�ǀH�ONONS)Ю������CAM_PAR�AM 1����
� 8
SONY� XC-56 2�34567890�Y �f�@����?�W�( С���8�h�х�ڎ��HR5ǃ��	���R570�B�Affފ������ڟ� ǟ�"���F�X�3�|����i���į!�CE__RIA_I����5��F��;�Я� ���GP 1]����s�����V�C󠸾�����CO�C ��(���ǀC8��@��H̺�CCX����Ch꺰p��x���� +C�����Ⱥ���+�=�G��ށ��HE>/pONFIG=�f��G_PRI 1�B�$r�����������(�~�CHKoPAUS�� 1���� ,wuj�|ߎ� �߲����������� 0�B�T�f�x����D�O���T���_MORGRP �2?� �\�� 	 �,��P�>� t�b���5�����eҒ.�?a�a�����K(���d�P�V��a�-`�/A�

s��������b&�i��ܦP�DB�����)
�mc:cpmidcbg��:��&�%y���p�U�   �  #�s*5� ���d܆�݆�ް{C�e�����{g�+/�/�{f/s/i��u/�
DEF ̋(K�)�b buf.txt�/�/���_MC������d,53����|ʇ�Cz  B��p�B�Z�B�X��B��~C� �Cޢ�D3��u
q�Dv��D�:�"Df��E�NNEA7E�V�ߓ=F�pg�F=C�Fi�W�G���Gp���G�3O�?L���
5����4P���N *B~��%�/��ʄ3@à1g/  TB�D�V@�a  EI�5� F*� F�G�$ˀF[� G�R�kNGl��G���G��&H���G֓�H��߃]��  >�33 �ށN�  n^��@߂#5Y�Ed��A���=�0<#�
 ��_�*2RSMOFS��.^�9�T1��DE ���l 
 Q�;��P  0_*_>T�EST�"__��R����#o^6C@A�KY��Qo2I��B��� �C�qR!�bT�pFPROG� %�S�o�gI��qRu����dKEY?_TBL  6���y� �	
��� !"#$%�&'()*+,-�./01��:;<=>?@ABC� �GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~����������������������������������������������������������������������������q�������������������������������������������������������������Eъ`L�CK�l���`�`ST�AT�c_AUT/O_DO��O��INDT_ENB�;���R�QY�K�T2����STO�~���TRL�`LETE��ފ_SCRE�EN j�kcsc 	�U�πMMENU 1�i  < �l�ol�K�u���FS ����柽�ϟ��� R�)�;�a���q���Я �����ݯ��N�%� 7���[�m�������ɿ �ٿ�8��!�n�E� W�}϶ύϟ������� "����1�j�A�Sߠ� w߉��߭߿������ �T�+�=��a�s�� ���������>�� '�M���]�o������� ������:#p�)+�_MANUAyLӏ��DBCOu��RIG�$�DBN_UMLIM�,1�e
�PXWOR/K 1k�_�-<_N`r�TB_�  m��Y0|�_AWAY�%�QG�@b=�P��_AL� =���Y�Ҁ��`�_�  1}!�[ , 

�:&d2/o/�&�M�t�IZP�@P�#OoNTIM��d���&�
�e#M?OTNEND�o$�RECORD 1�'kU2)?�!�O�?1-?&k�k?}?�? �?88�?�???�?c?O *O<O�?�?rO�?�OO �O�O�O�O�O_�O8_ �O\_n_�_�__�_%_ �_I_�_o"o4o�_Xo �_|o�_�o�o�o�oEo �oio�oBTfx �o��/��� ��>�)�7�t�� p u�����-��͏ۏ� ����N�`�Ϗ��o�� ��)�;������8� ��\�˟ݟ����;�Q� گI���m��4�F�X���TOLERE�NC�B�	"�L��Ͱ CS_CF�G ( +x'd�MC:\��L%04d.CSVY�� cֿx#A ��CH�z _/x.��G��},��RC_O_UT )�- �z/��SGN *���"��#��17-JUL-25 20:52���27-MA}Y��14:38��]� Z�t������x.����pa��m��PJP���k�VERSIO�N ��V�2.0.11~+E�FLOGIC 1�+� 	d���ٓ��p�PROG_ENB�2��WULS�' �p�_WRSTJN� ���"�EMO_O�PT_SL ?	��]�
 	Rg575x#?�74D�56E�7E�50i�dԂo�2E�d��j�"�TO  .����k�[V_� EX�d�%� �PATH A��A\��M�_��~+ICT�F��, '�`��eg��}�STBF_TTS�(�	��E��`���� MAU���ߧ"MSW��-D )��},t���.�!��]l�R�v������4SBL__FAULy�/�|�#GPMSK��^�"TDIA��0����`���!1�234567890xS�l�P��� ��//%/7/I/[/ m//�/�/�/�/�/LZ0PV �� �/�2?X?j?|? �?�?�?�?�?�?�?O�O0OBOTOfO8<x�U3MP$�I� �A�TR>�O�@PM�E���OY_TEM=P��È�3��4󜐰�DUNI	�w�Y�N_BRK 1���x�EMGDI_�STA	��GUNC�2_SCR 27[��_�_�_�_�& �_�_o o2or�nSUQ13y_+?|o�o�o�o�lRTd47[� Q��o�o���_>Pb t������� ��(�:�L�^�p��� ���� ?Ǐُ�0�,p ��+�=�O�a�s��� ������͟ߟ��� '�9�K�]�o������� ��ɯ�����#�5� G�Y�k�}�������ſ ׿�����1�C�U� g�yϋϝ�ׯ������ ��	��-�?�Q�c�u� �ߙ߽߫�������� �)�;�M�_�q��� �����������%� 7�I�[�m�������� ��������!3E W��{����� ��/ASe w������� //+/=/wa/s/�/ �/�/�/�/�/�/?? '?9?K?]?o?�?�?�? �?�?�?�?�?OK/5O GOYOkO}O�O�O�O�O �O�O�O__1_C_U_�g_y_�_�_�_�gETMODE 15'E�fa t�|�_GgRROR_PROG %�Z�%���HogTAB_LE  �[1O��o�o�o�ZRRSE�V_NUM �R?  ��Q�`�a_AUTO_ENB  u�SZdw_NO�a 6�[��Q�b  *�*6p�6p�6p�6p�`�+5pOastHI�S�cXa�P{_AL�M 17�[ �2��6|6`+t�@��&�8�J�x_�b.p  �[4q�R����PTCP_VE/R !�Z!6oZ��$EXTLOG_7REQ�v�y��SIZ�܄TOL�  XaDz�r��=#�
ނ_B�WDo�%��fQ���_�DI?� 8'E�t�TXa b[�ST�EPg�y��P��OP�_DO�v$v`F�EATURE �9'EQ��Q�Handling�Tool � D�ER Eng�lish Dictionary��7 (RAA� Vis"� Ma�ster���
�TE0�nalog� I/O��p1�
0�uto S�oftware �Updateb� �"/�k�matic Backup
��d
!��g�round Ed�itB�  25L�Camer�aT�FX� "Loμ�ellT��L,� P��omm9�syhۡ�h600��scou���uct���p�pane� D�IF���tyle selectѡ;- /�Con��9�?onitor���Hd�tr�Rel�iabT�ϣ(R-�Diagno�s��Q�	�H�Dua�l Check �Safety U�IFc�Enhan�ced Rob �Serv��q ��v	ԸUser� Fr���T_i��xt. DIO� f�fi�� )�\��endܰErrzu�L��  prנ�*�rO�� @���E�NFCTN /Menuİv�����.fd`�TP I�n?�faco�  �
E�G��p;�k Excذg�C���High-Spe�ܰSki��  P�ar+�H���mm�unic��onsn��\ap��urf��?�X�t\h8�U���connZ�2�Т !�Incr���str)�8��M�-6�KAREL Cmd. L���ua��}��B�Ru�n-Ti�EnvB�(<�@�I�<�+��]s��S/W�"H��Licens�e���� ad���o�gBook(Sy�>�m)	���"MACROs,�¿/Offse\�fĜ���H�!�Y�M1��MechSto?p ProtZ�3�o 5
�Mi4��Shif\��B6S�MixܰQ�����H�Mode S�witchY�MoTk���.�� ��Mt�Q�g�� �5��ulti-T�������)�Posj�Regyi>���  ! �}PA�t Fun1מ�6iB/��R�NCum�Y�3�G�P/�|�� Adju���	�/2HS�)� yo(�8�tatu����AD ��RDM�ޱot�scove&� #e�v�㱗���uest 86�7.��o�\���SNPX b��Y��Þ)�Libr%�
�r't I���� "���Ҫ�.S�o� ��s in VCCM����� j������㣀/I�� 71�0�TMILIB�X����g�Accܨ���C/2�TP�TX�� �Teln���Y@����K�PC�Unexce{ptܰmotn��� ������\m725����w�5����  h640S?P CSXC�i �� j*�� RIN��We���50,���vrl�زme�n" ��fiP-�a����P��Grid�{�play F �O/��? ��ELR�;�|�20��OR�DK�sciiw�l�oad�41d�s�t�Patd��C�ycT�h���ori�ɰ:�7c Data&� qu6�2�0�*�p������FRL�amc�K�HMI �De��(����k�P�C�φ�Passwword�644���Sp�����D#YELLOW BO�	�?1�Arc%�vi�su����#ti�OpX�^�! 2��aO��po�� t��ֶT11o�����HT���xy�	�   $�t۠ig��10�Ơ 41\+�JP�N ARCPSU� PR+�8b!O�L0Sup�2fi�l� �!��E@-�;�croc�82��v���n$ 12jSS0]e4�tex-� I��7�So��tf�ss�ag�� e��У�P���,��� "Tc VGirt��v�!�����dpn�
�J3ނSHADf0MO�VE T�MOS� O TԠg�et_var fails l�>PU�~1E���� Hol�d Bus %�h���VIS UPD�ATE IRTO?RCHMA A�{��vYWELDTV S� ]�DtS: R7[41��ouiPb}��y��BACKGR�OUND EDI�T "RC$REPT�CD CAN C�RASH FRV�R 62z1�SCr}a��s 2-D���r ) "��$F�NO NOT R�E��RED �` �m ��JO� Q�UICKaPOP �FLEN m41�S�Loc��gRTI�MQ%�#�FPLNs: FG��pl m��r`�MD DEV�ICE ASSE�RT WIT P�CV;PB�AN#aA�CCESS M �.pc��Jo��Q�ui±�Kbldm�gUSB$ ��t & remov��� Pg�SMB N�UL� ;a|�FIX���C��ACHIN�,QOL�`MO O�PT ՠa��PP�OST0�WDU �C�wQAdd�`aYd���0io�2��k$P�`W\0.$0`�O�IN&�P:f�ix CPMO-�046 issu5eC�J/aO-�0�r7130Т- ��vR�SET VARIABLES-P{��R�3D m��vie�w d��M��&�e�a���b��of �FD�5P:N@x �OS-1y0`�h isc���t��s t�3lo��7 WA�PZ��3 CNT0 T��/"�ImR�)�c�a �Pu��POT�:Whenapew�B�STY E�{1t���ptKQdo G�ET_�p �p��V�MGR LOl�REAd0C~QW�~1��(�l�s�gD�ECT�pLpING IMPR�DR(p+PB�PROGRAM�E�RIPE:STA�RTU� AIN-�;�ӠM/ASCIyIzPÂOF Lq��DPTTB: Nv�pML$me P����`:x�mo&�a�llW`!�ӤTorBc�A�U�HC�iLp�Ըth�`n�@ c�h��/GEA�!�toyu͐�RCal���k�Sign`� N�D�ԗThresh�123��`��09p : MSG_P��+0er  �Q�Aܠzeron��0� H85��RImlA�n�2D��rc�0�I��OMEa`�pO�NaP5�  נSRGEG:FF-Д� ]�|'���KANJI���n��J��c�0asn� d�!OA imm�c �INISITALIZATI�����~1wem����d}r+� LB A�U�Wqminim�r�ec[�c!�R���m>$�ro -1>ѮS�ܰir��@ұJ�1pdETw�� 5`?�I��ow u��< se� 1lc��YbPM ���p�Q���R`vR&��lu\�3�Re 0��4q�q1#���m <a�arn��ঁ?Box fo��*PORWRI�PW�S���v�09 F�pup~�de-rel2 �d�p� j��`━b�etwe��IND� Q���igE s�nap|�us��s�po TME��T�PD#�DO�p#aH�ANDL 1\kP�`vR��ȀD�ny��S�v�Yopera�bil� �T*�: IH � l\p��Vq�Hb�R�< p�a*�c&2�O�`FA,�.�-QV�7. f.v��G-T�pi�s��� �ɠtmLine-Remark ^�� RM-�` W��#SPATH SA�+PLOOS UIqFc�+5f fig�pGGLA����Vrp�������U�0ther|�V� Trac��"�tW�\b�s7��d��t�� n�@  ����3:���dK�y���it k8�d�P;ayR![2]�ü�1: g��s��d�ow�XQ��0IS��q�qEMCHK ?EXCE C���OMF +�Xah�� 35\k��)���QBt���'b���2[�c���e �`k�<�S�� BUGr�:�cD$`PETp����f�c4��0XPAwNSI��DIG���@OoPmetTCC�RG EN��CEOMENT�A M̀�K {�`H GU�NCHG �`� ECXT�P�2�bQS��93 wP8�x�OR�YLEAKq  �H5gyq�PLC �WRDN R �O9 /u�QSPE=p��G*�V ��$�t�n720\3pGRI��A�rT�PMC� ETH��pSU<7p�`  j5/n�/PENS�PN,���*P ont�`BR�OW�`!sRMV 7ADDz CN q�DC���PT3 A�LA2@ ���pSV�GN EARLY8�R��ŰH57�Ga�JLAYҀE 5(@M�PPD�p*@�H�S I`P�OGUCH8���V�F�q��comH�x ��E�RROR� DE �nJ��RO�CUSRS8pI��N4<q�-158n7�ORSR xP#aUp�P��Rqy�T�Fz��;�pk��t�� g�Ղ�B�SY RwUNN�  a�`��BRKCT�!RyO�p3@ \apS�Ƣ�AXxP���h8x+ q��ISSUrp} sPX�PTSI��K1M10_�IP�SAFETY Ck�ECK[��Á�������<#X�� �T�WD2�@�@�IN=V��D ZOp�5�X��t�DUALy� "M6�0�"r�F#�E��dPdNDEX F�t*UF�"Pʀ�0s�FRVO117 �A�PT6�KtqFA}LPTP2477D�6_�P�!;HIG�� CC�t;SNPX� MM��tq�d~�Vq�q#�
"��DETEC�Tq*@RRU�qA�P�5p
�9 y�)<9���7�T��Pds� �k�	���!Q����� t\4A�;A0�27 "Ke@" 8@HI��qXF8@4@H�PRDC"�
�aMB8@�IXF�b���zOX@8@����a�G}E�B�Ccsc�r�J8@�Ndctrld.�A�NZE�A5�I�Q��!�`�Df8@\�`m�878�Q-;� ��� rm`�
���PR̠78�@RaI8@0q�Q (~\�Mp��0t��!{B8@\PtQ<OX�St0�3hB�3nO�Vtp�A�@L�CF�L��� �Rplcf���J8@�WTa�mai�E8@mubov2_miTA�O�S8@U`�T[tT�AqPr674�xSShape G�en��8@j�I�[R��`�@8@T����%q 1(u8@��II�^�Q�~C�a�[8@;Ynrsg:0�4� � 4�CtMSr68@�r5hB5�z�Vnretsp "�r�Po�wng0bGCRE�Ka�ޠ��DAT�E�k�cr�eat.�q�M�a��oksqgtpadx1P��(�tputZj@�{�������܆28@`����Q����sl�ov��� �hexH��TB�8�ď�keyH�8@�pmZb�NR�1u7A+�nrgc8@UQ��pp�bUZ�dp0aj�921xSpl.Collأcq�\A��R1Nq�UA� (J�8@ip�_�WA��_�Y���a7hB7�ͦtp~[� "TCLS9o<Kb��clskyh[:��s�pkckZd� ��$�TQ���dA�rx��710a- KAR�EL Use S=p�FCTN9�a�a7l�0s0a�� (�� �a��~C8@��MI��c�8hB8"   ��8@ v	��v	   lomatea99�q�M����E�mcclm5�CLM;�� �j̕�E�et���aLM�	�h�yasp,���mc_mot�B�N��`8@H����Q��su'���Q�ȕ�䅮���jo�i#�ߕ��A_loqg�Z���trc�B����ve�ϓ�v��Q�WX��6�finde�rxSCenter� F1�lSw520���ha6rX� (<�r1,�Q�Ձfi�Q � NH0�I�ۡ���A8@uL���tq�a "FN�DRVϳ���etgwuid�UID�C 8@���������TA@�nuf;��P���ƞC�B��_z�Ӡo��q�G������l���fn�drTY��2䁴tcyp"�,qCP MF�:}38@517��6s38�E��gf6�� (��K��Q��-�X��A&�tm6�P�İ ��Q���	�͘���tm�Ĵ�b8@e0j��TAiex��aP��Aa�ذ�cprm�A��l�_vars��
��dwc7 TS0��/�6��ma7AF��Group| sk� Exchang�J 8@�VMASK �H5�0H593 MH0aH5@� 6� +58�!9�!8\�!%4�!2���"(�/�@�;OMI� `@a0hB�0�ՁU4U1#SK (x2�Q�0I�h��)��mq�bWzR�DisplayImQ@QvJ40�Q8aJ�!(P��;� 0a��0�Ϙ� 40;�qvl "DQVL�D쌞�qvBXa`�uGHq��OsC��avrdq8�O�xEsim�K40FsJst]��uDdX@TRgOyB�Bv40)�wA�~���E�Easy �Normal U?til(in�K�11 J553m��0b2v�Q(lV40xU)���������k98�6#8Uϕ�|�rP "NOR��dw d.a}oKksu�O�W���O�Y�W`�j0�6�H� mOenuuyP6�M�`�wRX�R577V�9{0 �RJ989}��49b\�`(�fity�����e�<?L��Vsmh`��8�� C0�Sv�q�8����w�pn "MHMN<��ޣx�Ay`�o�3@�u�`f�І�x�t���tRzQ��LV��vP�tm���|I�1{oPx ��2|���I�3I/B�ogdstǏًmn吼���}ensu_�L<���h!!��Rt��?huserp��0���ʐcM�_l�xP�oxe��рpoper��|��xdetbo/� l>�x���Ps$p�`����OPydspweAb͓��z'R��u�Rr101&S՟{t�`12�Z4�30���D���`4�
�4�5���KQ�m[T��dUCal G40`�Q)p40}������9;��DA��� v	LATAu�mpd�\bbk9�68��68c�fb\l�41969y�9�|��D���bd� "B�BOXêM��sc�hed����m�se�tuM:�����ff ���40��n�41�ϒ�40q�col��|�1�cxc�ؘ���li�� X�0���j��&�8�4 �<�ro5�TP E��#��ryK42�r��;�(T+Q �Rec'�ʈ1Iw�84������Ak971���71�;���parecjo��QNS��[T���dXrai=l| nagek�M �,QT2 *� (�ĜR%<x�80!�bh��p��4��4��yDgl�paxrm?r "XRM�g�l�brf{���n����kl��9turbs�p��㧑- �l0195	�g�625C�M h�+���)89��	+��B6��o�ҹ���x�7�q40����pd "TSPD�=<��tsgl��l��:dQ���8Bct���K�vrE�aܮ�����  c�!���21�`�( AAVM l�2�0 �@fd �TUP him �(J545 �l)�`8 616 �%�VCAM ���CLIO �(�0:�5&  {(F\ MSC �R�t"PBsSTY9L�D!28 :2\ �NRE F2h SC�H6pDCS�U tpsh ?ORSR �rD!�04�SEIO�C& \fxh 54�2 LEX"� E�SETn�8!H ��s�h8 7H �M'ASK�Ø"7>���OCO*`x�!03P"6�!/400:66$ �G639.6[8LCH�!6OPLGR703�
5MHCR��0CЄ (! �06�A.f�8!54
��00DSWb 588�180 ��h!37 88 (%D�"02C24���2'7 q9�25��2�-6�05��9P�RST bBFRDMES�!zB��930 _ NB�A  6� HLBo 3 (~!SM�@� Con� SPV3C �8!20z���TCP aram�\TMIL �A��@PACETP�TX �@p TE�LN 96��29^�%UECK��r UFRM et��P!OR ORP IP�L%CSXC�0j��1CVVF l �FQHTTP satA")�I#� CGHP�8ZIGUI��0�hPPGS T�ool� H8�@d�jZ��!@�h!63��%�@32Q\�31 �B�h!96�%R65�1�Rs�!53 T7FAD�R41�8"[1 ��oo�"9��41775�"/@�P�VCTO�@�U�!s�h!80�%PRXY<�R�!770 �b8 ?885 ol3P� L� аdi� �`ڳ�h LCP{Q� TSS �b�26:����@�CPE �HT@V�RC~�tQNL <��@002 %��b�	0dis� �`7 `<��a\0�T�`1 �`{en�b4 652�`)FU02Q0Πo`dp�Ptu�r4 $�r5N��RU0p@n�se�QJp1 AP�FI[ Jp3�g34>�g40 alxrlE1t44w46� ts U0  7v�0�O��r5�e�p7 po "sw�a61:���r4��r5 QpwGr`�$�p8R�"sP`�tQ�b�36w77��w8`�v83���r8��&:��pOq8�8 "/rkey8�9F��a;90�91 p�#@���� �D095�g9-7*pur�A1@d����P|P�q1�0Qpl�Sq1p#4��]a!s1&@sl༂8�Ӽ�$\1�d1�`��v�@�{�14p�ae��5 �h2��`�6ޣ��7�f1p@��d�YpCqd�ـd�1�`uq��� BCu1< Oq� ��7ReU1$ �u1�Pϱ� ܺ�@- WQ158 ase C���9 B��60 8�2ń�p���4 (Wai��`吢!��i7E��8�EU1P`�ro9�<�1��<�2 ��<�	0��T��l��5J�l��cC���9�%�MCR��P�2��`�Q2@967��Q��8��9Z�2�TPB���P�2P7UA5@�o���
�5�`U���3 w���?AH�E�1��c�qAwl���A�1��512 f��1�u5Р���a5p$��56�+a��bQ5h��Ұ�1 @���pp�b[�538� xaB��|p�4�2��11/q5�p�4U5�P16 (߲�Pz��0��8�P����$�p�e5`�e5(�/�P`bbf>�X��$Z��U�5d�\� ~X�7 	  �ÿ8 k_kv��7s9 s�82 &�H5��E6���p����Ah���ñ���3J"ܫ`��4 3Ȥ59Jѧ6�0t���8��q6D0$�$�4 7���!���<�j670\tchk<�Ps0��<�B<�90��7�H<���<�\K�<�q�� ��A�C<���q�<����<�t��sg<�lc$���FA<�H��<�`��<Я���<�hk�� <Щ�B<е�o�<����<��K�<�dflr0��<Ш��� ��oҠ`���D�;�<�gEvam����B<г�o������<а�KЀ�creexl����P��<���|���j6<�s��prs.`���\���<�7������f�sgn��P�b�t�at��<�L��1B >!�svsch/  �Servo S���ule>�SVS��44�1u�_<���� (����ched���,��~��A\�� �� B���B�qA�����cj�� � 5��1<���Ә�p�css "ACS<� &(��6� �����c el���Q���~��torchms�n<�- T�Ma`�x����09 J5;�598 J681
s�7� 8��b���<Чa����te,�s�����/�E��s m��ARC.�� 1q�4�!=��C�tc�pA�@t�L��f� F����7#�2x�SE�r����UtmS�0960'���RC���`���� p��96G0= '��"H5W�� ��L���\f��� �PATb���`!40U�#!Stmt��E ��� �pMA��!p��z�2?�inA_<�X��r�X e/	cW����V���чetdl�vߏ\oveto���܏��mmonitr�0\��|#�0st��?.6a��PP����! Q�!y`�`am9e �Arol�c�43�0 �p��6��01� 25��  �<� ?v	�v	�A@�818\n; <s��I�B�2�pMPTP�"��C�1mocol��,��CT�v�'!� 0�A���8P53��y`_Touchs�s�`��<��J5���� �`mP����n[PQ �a,�E�a��IP&
&�Pth�A<�KF#R��m;�Qetth�TGHSR'�q-�Rt��o "PGIO�#�!$s�ISwka�"W�K��!�MHqH+54��5w5n/�Sm/��@ 7�*�da���8`!w/Ac��tsnf Tk�/�#gb��a��u`��^m�`u ��Zӭ�ܱQp�є� #���Ka<��M��t5QtZ�a<��dFS�5GK����G�1or��dW��64��tPx� ��P ����x,�� ?$���P<�Z4e7�g "SVGN.o�x�copy "C�O;�Wj$�O�A�9� "FSG�ѧ�%7���_��f� wQSW�F*!"(�sgatu`ɀ���_
��tp_�TPDo��9�7�9�#dߎ?���h�G�AT���!#��  �Гf�` ��" /� �w�Z� �b?6?�  ����� ���E ���M� �chrT� �K6K� �sms� �o6��~��gtdmen?3� �?��� ���mkpdtd2 ���, ���pdQ�X� ����� ����mvbkup.� �[�C�С��mku�no��prp���m�kl �4��s �n�iU��� �ldvrw���glg�4�� �p�棑��aut7�.pб�旐 �ַ������su3� �Ǜ�  �Ƿ� ���\ �6�b2X� ��&�� ���<��A4�  ��B�   946"� ��fB� �t\pa�ic\p4k94�7 ���F#���� �i�ctas���pa`���cc:�<��o������gen�� � $��F�lnp � �����stf@��1��wb�O�c��Ջ�`��߄�vri�ߢ�а�-T�� ���p�flowl� OPAc��ow���R50qtS �#T� (A��4�#���pѣV�cu3�QF�� ��SI�ac����4�6����s&��pa���!!���� ���55 �b �o)�p���0娿>
�afcal3�P߁ ��f��}���`�f��m	߳�p�d�m�/���a/��$C`ѷ��� �! track�\P� 0�ine/R?ail Tr�]T�J�69W�T  (L ��8(`љT.�`�%���D��P0� (��8�48��_ɛ�⇒A4����� �3�b13���alV@ ��NTf���%��Ii�n]0m���aen ������&?5�c@Itst3@��$� ���`�,R9�%����0氱%��pop_eners-OW �dDev��F�M�6 W���|A�Pc"�l!esv� �,��R��V$��Q���U<�V$ �k9j �6��# ������%paop/!OP�NU�V ��2celL��8g_��/�6��tscG��$���V!�3� 5vro!p�ߡ�7`�n(`� V"2D�a V'O$:S|9��� PumpE� �jQ�@�" ��!
��@бMSC#�@��)P��A�C�`��� � �v���� \mhplug�@g�"7Pb��uK")㠱io7��CJ0��E�LIOj q1g 7A93շ��5 q9 t����4.rb ST��R��CP�J989�P�LSQE�' �e C3Q(P �/Ov���o�P�� ? I1�R���5�5��f�I1`�tcm;io��MIO������Utco1"CL0�1V �cBK`io"��uM?���Sl�I0�ߢ�Eg �o���f �1tI4\onfdtI����e%�p27�Int�e�TB CoMo�o1E�R�(do5�54 (;r>Ex,p��nR##ipc�/L>��qp5���
oQ é�1�p����7/o��j�ra�pd�CDV�_��rP�֮��qp2c�nd��s �p��a �o�r`҄�S��"�c�1a�c���2kIԿ?A�pcrt���or0�qd#��"���3p+�཈D��Џ��vr2k�0���AG�.+�η�cho�;�uCp��(� �uV630� fwe P�mී�@���,`��TX�� ��d�chp "_��(	�3�����8����\p3�v����ш�9�3�1 ������low�[ͧ���chk���㳦s��s?Ө0�i�1h���2��i�w����s?1*�-0	�:�O��vr����৓0�'���PFRA�PWat?1rne@E�P�sp�& ac5� \_A�rbo#�,�a ��g��������Q=s<�ICSP+ �9_����� �q�F�A9PH51IQK93 7��HX6hQ�]PVR`S5��fPR6� iQWPR� (P^!am S�u�"��A�I0�tpprg��0���`h�@2atk932�!��E�^�^�asc "8�C��S>i�atp�"�d��@1I�
g�dsb�lfltJA�Qsable Fau�P{C!��EV0ex/!?DSB (DC��t�$�p��X 7�  �� 5��Q�t3*�~l���td9� "!0%�(5��sb9኏���\	�6#���@5��p$D@550-Ad�just PointO"tVJ�Rs�z�@䐄��!�X_�Yj�^�0\sg��4�߼}7y�\ada�"�ADJ���j�Qe�tsha<�SHAqP�sŭ'jpo�r 4�t�!��$ ��C�|�	Tk!bRPK�AR/Qiagno�stì!O!vV6�6 J`ew0�(��L���/�&krlde� ��PP���h�U b���r3�Pp<?q��DBG2C��� �X�o�1U��� ��WT`�@ip�JCM�aipper� Opv`1Se}78 (MH GF�  ;":�&##�� a�xX�֕$��388C�P����#��9.�9C�H�g##PPk�Q��8�! �_"$�"��=0%�P��A  $��_�#%0AQ�C~2� Mat.Han�dlE��!= &�pq MPLGET�0�1(�3�Tt&P�Sٰ'�B �1��B0����&p��H ��PP �'p��@�C7�PP	�TG�tD5�}m��q�Afhnd "�F_R  ���|��PP	   xT�?Q���P(Pa��TAo�����?�pmp�aO��JP ak92�5��2`@O�JRp�sQ`B2�unLHP�Tgse�GSo1�O�W�QT��v !�R�P�tp~���JRdmoan.�@��V�!ns�hYvr�QJ�g�Q�o��jY�HS~7sl�f .��pen�PDnR(R8&���ɐ823'�� ٔq���g� ���� 1��� S�� ? �c\sltQ�!|QE�P��a�r�tPg��P�� �v��"SEDG8�s0�qtdgY T��� �vP`ho�s`<`����qc�`g
�e` op�w�a@o"�ile6�H�e�ȅnR�� x�e! j517�>Ճ��J%��e�`��Q4��Q&�L�!F�J�=�o�5�z/l17���_�œ���`C0C�  ���LANG j��A���8�����gad��X�#�jp�.�0�4�Ē�ib���s�Ƒpa����&���j539.f��,Ru� Env
������3H�z�J9�����@h�Ф
Ҕ���2�a2���� (KL�n-TimФ�⠤���p�3�TS����\�kl�UTIL"�o���x�r "QM�Gl��!������1� "��S�T3�\kcmno��SФT2����ut�.�lrgeadc�}�exY�(ܤ�r��\��l��Ф�w�3��2C�*� - �C�D�E!Ĥ� .��C� R CV̴�Ҁ�C\p�Р���pďtbox��.�@�c�ycsL�:�RBT�E�veriOPTNE���;ӕ�k��e�ߦ�a�ߦ�hg��ߥ�DPN��gp�.v��r�ptl�it��0�4��te\cy����tmnu3`�r�����5UPDT��������駣��i�te �� swt�o�,���oolB �F"�Y���Q��(q��gr3��䪒��"�䴁w������߳��s��������������lS���bx " O�� ����l����0P���A�l\t�� ���������	�Colr�e!��R C��r��&r �m;`��Chang�Lq�T1 �rcm3�"��
�� 6���"����sP70���"��22!2��2D4�57�� CCF�M�H��accd	a��Q�c' ��K�@�0���K!����mo! ���,$Á��!"
 ����/�/����	Y�`,$��)�,$sk����m rC%tS1,$+�x��k1�%unc.,$poñ�1��sub��p����1��cce�5 /!&��-/?-W/i&vs�}/�%#�#�/�.@C��/� C%
�@? U ��&+��F:qt�
pD�Ѓ D	 � U�:7�Dxmov.�P��DPvc5Q.�tfr@PeC_UY?geobdtg_y[�tu���P���PTUt$�P�Sx�_�^z�_�\gvar�_�\xy�_.�[pcl`c�P���P�Ue�Pgripssuaoskuti��|�ovfinfpo}��o�j�b�P���Qud�\�aX��Pc�\Rrp��Qnƅ�P�v�P)tm�#qƆ�P�v�a+rog��a��\Q�?a+rpal?a{�{spa���P �u�Q�t�_TZp�0�osipkag3r�ovlclay(�:�t�pT�d�pu?a�c�A������KtKa�P��r��qTf|rdm���{rin#r���s � �2���|s�Pd�&v�tv��v�h�0���ystn* џ�yt'�1�p��D�p�uϑ�#�ul�@o�W6�2�siupdl�]�o�#vr�on��`1L�zp�`\�r���il3F$|l4��ǉ#q54�FyB�Տg{�`���{w�cmס���wxfe�r�UYtlk2pyp߿UYconv���sicnv�Qʯxaqg��H�Z�lct`a�o�=�p��׭nit�0믁�3������ � �� v�	�v	$��a�lϑpm�r&�B�e Wa���f�%���� ��I��߬�u�ͬ�Ka�mT�f���c��w��roǁ#�5�����?� sm��y�a��y넑 ������`����͐ϑ��p��m�Wa�1� ��A�6�S�e�X��� ��\Q}����������� ĥw߉�西߭���� ��#q0��rs�ew�@��1�a��z긱n@��.�۲;�d�������  � A�d	T$�1 pc! P��e �e� 	lf@C�@��s/�  ?�����8�� �������re�g.�C=��o�99 ~@�����$FEAT_INDEX  z ��e�� ILECOM�P :���1!!z$#�SETUP2 �;1%;"� � N f!$#_AP2BCK 1<1)?  �)��/��/  %�/�/e 4 �/�/>%�/$?�/H? �/U?~??�?1?�?�? g?�?�? O2O�?VO�? zO�OO�O?O�OcO�O 
_�O._�OR_d_�O�_ _�_�_M_�_q_oo �_<o�_`o�_mo�o%o �oIo�o�oo�o8 J�on�o��3� W�{�"��F�� j�|����/�ď֏e� �����0���T��x� �����=�ҟa���� ��,���P�b�񟆯� ����K��o����� :�ɯ^�����#��� G�ܿ�}�ϡ�6�H� ׿l�����ϝ���@)�t Px/ 2� �*.VR��߅�*�@߂�F�j�T���PCrߛ߅�FR6:����V���z�T �!���K� x��q�S�*.F�D���	�Ӑ���^�<���STM ���'���S���i�Pendant �PanelS���H I���9���U�������GIF0;���8�����JPG���;��]oR�
A�RGNAME.D)Ty�>�\"���Rc	PA�NEL1Y�%@>��e�w��2��A/�//���/�3 _/�/��/p/�/?�4�/I?�7?�/?�?�TPEINS.gXML�?>:\�?�t?�1Custom� Toolbar��?Q�PASSW�ORDg?w�FR�S:\:O�? %�Password Config{O R��OSO�O�O��_�O B_T_�Ox__�_�_=_ �_a_�_�_�_,o�_Po �_Io�oo�o9o�o�o oo�o(:�o^�o �#�G�k� ��6��Z�l���� ���ƏU��y���� ��D�ӏh���a���-� Q���������@� R��v����)�;�Я _������*���N�ݯ r������7�̿޿m� ϑ�&ϵ�ǿ\�뿀� �y϶�E���i���� ��4���X�j��ώ�� ��A�S���w���� B���f��ߊ��+��� O���������>��� ��t����'�����]� ����(��L��p ��5�Yk  �$�Z�~ ��C�g�/� 2/�V/���//�/ ?/�/�/u/
?�/.?@? �/d?�/�?�?)?�?M? �?q?�?O�?<O�?5O rOO�O%O�O�O[O�O O_&_�OJ_�On_�O _�_3_�_W_�_�_�_ "o�_FoXo�_|oo�o��o�`�$FILE�_DGBCK 1�<���`��� ( ��)
SUMMAR�Y.DG�oblM�D:�o*n`D�iag Summ�ary+8j
CONSLOG q�n�=qConsole log��7kpMEMCH�ECK��2���qMemory �Data3�;g� �{)�HADO�W(�����C�S�hadow Ch�anges���c-���)	FTP������=��qm�ment TBD�;�;g0<�)ETHERNET0��`n�q~���=qEthernet �p�figurati�on��B`%�DCSVRF/��'�@�C��%� verify allC�ޑc1p� �DI�FF8��0�ůD�{%Z�diffǯ{��q�1������J�� X�q�|�	�CHGD�&�8��ͿD�ܯ�����2pĿ����R� `�yτ�GD�.�@����D�����FY3p�ϳ���Z� h��ߌ�GD$�6�H����D�����UP?DATES.$�
�~ckFRS:\"��c�>qUpdates Listc��`{PSRBWLD'.CM��blN���e��pPS_ROBOWEL\�6o+�=� loa��o����&���J� ��n�����9��J o���"��X� |#�G�k� d�0�T��� /�C/U/�y//�/ �/>/�/b/�/�/�/-? �/Q?�/b?�??�?:? �?�?p?O�?)O;O�? _O�?�OO|O�OHO�O lO�O_�O7_�O[_m_ �O�_ _�_�_V_�_z_ o�_oEo�_io�_zo �o.o�oRo�o�o�o �oAS�ow�* ��`���+�� O��s������8�͏ ߏn����'��� �]� 쏁������F�۟j� �����5�ğY�k��� �����B����x������C�үg�v��$�FILE_N�PR�]���Y�������MDONLY 1<��~U� 
 �� ۿ(���L��5���Y� �}Ϗ�ϳ�B����� x�ߜ�1�C���g��� ��ߘ���P���t�	� ��?���c�u��� (����^������� $�M���q� �����6� ��Z�����%��I [���2��~��VISBCK��|��ų*.VD�|*� FR:\�V� Visi�on VD fileVd���� ���	/./�R/� v/�//�/;/�/_/q/ ?�/*?<?�/`?�/�? ?�?�?I?�?m?OO �?8O�?\O�?�?�O!O �O�O�O�O{O_�O!_ F_�Oj_�O�_�_/_�_�S_�_w_�_o~�MR_GRP 1=���LeC4  ;B�`	 ��lo�~li`۬B���D��fn�ӺMT� �?�� ����e`i `a�o�khb�h�o�d�cic.OLp��L)I�K�w��M���HW'�E��|�i`�?�=tB����A��>���B(6�9���l}Aƌ�A����A��KA��_9A����p�l}F@ �qhq�y�~�g�fF6�D��MqD�� BT��@��Ô~xpD��6���l����5��5��|��~e9��B �B��A�.�BWqr�B�~�~-G*�A��B{��A���BI�$B�l叐�A�����A�܏e��P���t�  @��0@�� =(��@ܙG����� Ο��+��O�:�_����p�����eBH` �ā����8ү��'�d
���Z��WZ�a/�FX
�A@�~��@�33@���'�\��[���ѿ��@��񿋯�*���N�9�r�]ϖρ�<��G�=�<��m]<�+=~��m<c^��8�eN7��7�ѷ7�x7;��51���	ߤϨ�?߾d2^`Yb`�*b`�����F�`�Y�b`��B�0�����C�^o�߂o�o �߸o��o�� ]�(� ��l���������� ��#��G�2�k�V�{� �������������� 1 ��-�) �������0 T?xc��� ����/')�'/ M/_/q/8��/�//�/ �/�/�/?#?
?G?2? k?V?�?z?�?�?�?�? �?O�?1OOUO@ORO �OvO�O�O�O�O��_ ��J����`_*�_N� �_�O�_�_�_�_oo 'oMo8oqo\o�o�o�o �o�o�o�o�o7" [Fjh�x� t��!��E�0�B� {�f�����Ï���ҏ ����A�,�e�,/�� �������/�J��� �=�$�a�H�Z����� ����߯ʯ���9� $�]�H���l�����ɿ ��ƿ���#��O�OV�  _z�D_V_��z_�Ϟ_ ���
�C�.�g�R� ��vߛ��߬�����	� ��-��Q�<�N��r� ���������)� �M�8�q�\������� ����������7" [Fk�|�|�� ��֟3�WB g�t����� /�///S/>/w/b/ �/�/�/�/�/�/�/? ?=?(?:?s?:�LϦ? p��?�Ϧ� O��$O�� T?]OHOZO�O~O�O�O �O�O�O�O_5_ _Y_ D_}_h_�_�_�_�_�_ �_�_o��@o
�go*o wo�o�o�o�o�o�o	 �o-*cN�r �������)� ;�M��������� ˏݏď��%��I� 4�F��j�����ǟ�� �֟��!��E�0�i� T���x���ï�?�?�� O��?OO�t�>O ������ѿ��ο�� +��O�:�s�^σϩ� ���ϸ������ �9� $�6�o�6o��Zo��R� ���������5� �Y� D�}�h�������� �����
�C�U��y� ����d�����:����� +Q8u`� ������ ;&_Jo��� ���//گ4/�� x�j/4��/X�n/|��/ ��/�/!??E?0?B? {?f?�?�?�?�?�?�? �?OOAO,OeOPO�O tO�O�O���O�O_�O +__O_:___�_p_�_ �_�_�_�_�_o oo Ko6oooZo�oZ��o�o �o�o��xo
G2 kR������ ���1��.�g�R� ��v�����ӏ���	� �-��Q�/*/��N/ ��r/�/ޟ�/��/)� D�M�8�q�\������� �����گ���7�"� [�F�k���|�����ٿ Ŀ���O�O�O��W�B� {�fϟϊ��Ϯ����� ����A�,�e�P߉� t߆߿ߪ��ߪo�� +�=�a��߅�p�� ���������� �9� $�]�H���l������� ��������#G2�W}h�p��$F�NO ������W
F0� �  #��1 D|�� R�M_CHKTYP�  � �q�� k�� ��OM� �_MIN� m���}�  X� �SSB_CFG �>� ~�Jl�Aj|��TP_DEF__OW  m��>�IRCOM� ���$GENOVRoD_DO���n�THR d��d�_ENB� ��RAVC_G�RP 1?3� X�e/��/�/�/ �/�/�/�/�/? ?=? $?6?s?Z?�?~?�?�? �?�?�?O'OOKO2O oO�OhO�O�O�O�O�O\�O�ROU? E�. q����>��8�?#�O_�_K_m_o_ꐖ  D3���_E�_q�@A��\Bȡ��R���>Y_6 SMT<#F�C-�Ufoxo�o�HoOSTC,1GYn?��_ 	�hM�k�o�f�oyeCUgy �z1�������p	anonymous�5�G�Y�k� w��o�o�o���� ��*�<��`�r��� ����ˏ	����� &�8������������� �ȯگ���M��4� F�X�j�����ݟ��Ŀ ֿ���I�[�m�ρ� fϵ��ϜϮ�����}� ����,�O�Pߟ�t� �ߘߪ߼���/�A� C�(�w�L�^�p��� �ϸ����������a� 6�H�Z�l�~������� ����9� 2D V��z������ #��
.@���� ����������� //g</N/`/r/�/ ����/�/�/?Q cu��/[?��?�? �?�?�?)/�?O"O4O FOi?�/�/�O�O�O�O�9m�aENT 1H�[ P!^O_  `_?_._c_ &_�_J_�_n_�_�_�_ o�_)o�_Mooqo4o �oXojo�o�o�o�o �o7�om0�T �x�����3� �W��{�>���b��� Տ���������A�� e�(�:���^���������QUICC0 �̟ޟ?��1@��.����2��l�~�߯�!ROUTER�௼�ί/�!PC�JOG0��!�192.168.�0.10	��GNA�ME !�J!�ROBOT���NS_CFG 1G�I� �A�uto-star�ted/4FTP:?�Q?SOBχ?f� xϊϜϮ��?������ �+�߿�P�b�t߆� ��6�����(�J�  �1�C�U�g�6ߋ�� ��������x�	��-� ?�Q�c� ?2?D?���� �����)��M _q����:�� �%t�����m ��������� �!/3/E/W/z{// �/�/�/�/�/6HZ  ?n/S?�w?�?�?�? �?�/�?�?OO<?=O �?aOsO�O�O�O�/
? ?.?0O_d?9_K_]_ o_�_PO�_�_�_�_�O �_�_#o5oGoYoko�O �O�O�O�_�o&_�o 1Cogy�� ��oT��	��-� |o�o�o�o����o�� Ϗ����)�;�M� _�q��������˟ݟ��ÿT_ERR �I�����PDU�SIZ  �^ڴ��$�>=�WR�D ?޵w�� � guest+�}�������ů�ׯ��SCD_GR�OUP 2J�� �`�1��!怒L_���  ���!�	 i-	��E���Q�E� EATSWIL�IBk�+��ST 4�@���1��L�FRS:�аTTP_AUT�H 1K�<!iPendan�������!K?AREL:*���	�KC�.�@���VISION �SET���u���! �ϣ��������	�߀P�'�9߆�]�o޽�C�TRL L���؃�
��F�FF9E3��u����DEFAULT���FANUC� Web Server��
��e�w� ��j�|��������WR_CONFI�G MY��X����IDL_�CPU_PC�惑B�x�6��BH��MIN'��;�GNR_IO�K����"��NPT_SI�M_DOl�v�T�PMODNTOL�l� ��_PRTY���6��OLNK 1N�ذ�� �2DVh��MASKTEk�s�w�Oñ�O_CFG��	U�O����CYCL�E���_ASG� 1O��ձ
  j+=Oas�� �����//r.�NUMJ� �J�� IPCH�x��RTRY_CN��n� ��SCRN_�UPDJ����$� �� �P�A��/����$J23_�DSP_EN~���p�� OBPROqC�#���	JOG��1Q� @��d?8�?� +S?� /?)3POSRE�?y�KANJI_B� Kl��3��#R������5�?�5CL_�LF�;"^/�0EYL_OGGIN� q���K1$��$LA�NGUAGE ,X�6�� vA��LG�"S�߀���J��x��i��@<𭬄�'0u8������MC:\RS?CH\00\��S@�N_DISP �T�t�w�K�I��L�OC��-�DzU�=�#�J�8@BOOK U	L0��d���d�d��PXY�_�_ �_�_�_ nmh%i��	kU�Yr�Uho�zoLRG_BUFF� 1V��|o2 s��o�R���oq��o�o #,YPb�� ���������(�U��D/0DCS �Xu] =��� "lao����ˏݏ�3�n�IO 1Y	# �/,����,�<� N�`�t���������̟ ޟ���&�8�L�\� n���������ȯܯ�}Ee�TM  [d�(�:�L�^�p��� ������ʿܿ� �� $�6�H�Z�l�~ϐϢϜ�d�SEV� ].�TYP�$��0�)߄m�1RSK�!O|�c�"FL 1Z�� ����߯�����0����	�:�TP5@����A]NGNA�M�$�E��k�UPSF PGI|%�1�%x��_LOAD0G �%Z%TES�T_Z��MAXUALRM;'�I( ��~���#� V�#a
��CQ[x�8��n���"�1060\	 �F�	�Ϣ��������� ���� D'9z e������� �R=va� �������*/ /N/9/r/�/g/�/�/ �/�/�/?�/&??J? \???�?k?�?�?�?�? �?�?�?"O4OOXOCO |O_OqO�O�O�O�O�O _�O0__T_7_I_�_ u_�_�_�_�_�_o�_�,o��D_LDXD�ISAc���ME�MO_AP]�E {?��
 � 5i�o�o�o�o�o�o�o���ISC 1]�� �oTd�� \no����� ����I�4�m�� f���$��������� !��E�ƏT�f�:��� ��ß�����z��ܟ A�,�e�w�^������ ~������ �=��� L�^�2���������߿ �r� �Կ9�$�]�o��(t_MSTR �^�͂�SCD 1_xm�W���S����� ��=�(�:�s�^ߗ� �߻ߦ�������� � 9�$�]�H��l��� ����������#��G� 2�W�}�h��������� ������
C.g R�v����� 	�-Q<u` r������/ /'/M/8/q/\/�/�/�/�/�/s�MKCF/G `���/�¿LTARM_2a��2 ��#\`Y>G`METP�UT`�"����N�DSP_CMNT�s506�5�� b���>�"1�?�4�5_POSCF�7�>�PRPM�?�8PS�TOL 1c2}4=@p<#�
aA�! aEqOG]OO�O�O�O �O�O_�O�OA_#_5_ w_Y_k_�_�_�_�_�Q��1SING_CH�K  +O$MODAQ73d
?�7:~eDEV 	���	MC:MlHS�IZEs0���eT�ASK %��%�$1234567�89 �o�egTR�IG 1e�� �l��%��?  ` A$�ÜfYP�a�,u��cEM_I�NF 1f>7� `)AT&FV0E0N��})�qE0V1�&A3&B1&D�2&S0&C1S�0=�})ATZ�� �H�E��q9m��xAu���X�������� ����� �v�)���я��П�� �����*��N��� ��7�I�[�̯ן��� 9�&���\����g� ����i�ڿ������ï 4��XϏ�iώ�A��� m�������߿�ѿB� ���ϊߜ�O����� �ߟߩ����>�%�b� t�'ߘ�K�]�o߁��� ���(�_�L���p�+�����������.ONIwTOR�0G ?ak�   	EX�EC1�#23�45�`7*89�#�� xxx*x6 xBxNxZxf�xrx22�2��2�2�2�2��2�2�2�3�3�3aR_�GRP_SV 1�g�y�a(�Q����^?3>ӿ�^�l;�]�?�p�"�(;vHm�a_�Di�n�!PL_N�AME !�5�
 �!Defa�ult Pers�onality �(from FD�) �$RR2� �1h)deX)dsh�
!�1X d�/ d/v/�/�/�/�/�/�/ �/??*?<?N?`?r?@�?�?�?�?�?�82S/ �?O O2ODOVOhOzO�O�Ob<�?�O�O�O �O_"_4_F_X_j_|_t�_LhR� 1m)�9`\b0 ��_pb�Q @D��  �Q?��S�Q?�`�QaAI�E�z  a@og;��	l�R	 0�`4b@4c.a�P��Jd�Jd�Ki��K�J����J��J�4�J~��jEa�o-aƸ@��o�l�@��z�b�f�@��S��a�Q�o�c�=��N��
������T;f��
���m��*  �p  �$p�> p�$p��o?���?�����=����o�Bntr�Q�skse�}��l�p�  ��pu`j  �#p��vks��� 	'� � ��I� � � ���}:����6�È=���N��b@^�d��n�Q���{�R�x���nyN. ��  '����a�`@a�@�t�@p@p�n�-CpC0�f0�+p�B/pC3}�P��@%�Eab��oo$|m�/���gA%���. ���z�`�P���QDe���˟��(���m�� �t� O� ru� �4 �xR�c��s� :	e�a�P�` �?��ffb�!�����7� ��گ쬛af���>搠���iP��P;�e�S�Ea4f�u��>LX��s�b<	��I<g�<#��
<2��<D?��<��
vo���¯�S��S.���?offf?u�?&�ޗd@T���?��`?Uȩ?X����Z���T:z �TB��Wa�з*dů�� �Ϻϥ��������&�`8�#�\�h�+�F.  Kߘ�G߼�3���Wɯ����G�@ G����X�C�|�g�y� ���������jZ�� �ￏQ����ߙ��� ��3�������/ A��t_�����������b�� �@+Fp�IP(�t��%���[`B�0����<ze�cb!@I��
�M`B@���@`�9@y���?�h� ��@�3�[N���N�N�E��<��/:/L �>���ڟ�A�p��C�F@�S��b/DpX������@�t��%��h��`/qG���GknF&��FצpE,8�{�/ F�Z�G���F�n�E�DE,ڏ��/� ���G���F7��F��ED��.��C?.? g?R?d?�?�?�?�?�? �?	O�?O?O*OcONO �OrO�O�O�O�O�O_ �O)__M_8_q_\_�_ �_�_�_�_�_�_o�_ 7o"o4omoXo�o|o�o �o�o�o�o�o3 WB{f���� �����A�,�Q� w�b����������Ώ ���=�(�a�L����p�����(r!3�j�i��r���ꕢ�3�Ա�ڟ�u�4 ����u�Pq�2�D�&�jb^��p�1w���������ʯ���ܯ�� �s�P^�PD�c� `�m���y�\������Ӱ�¿Կ����� .�G����}ϳϡ� ��홍�U�_�J���$�y.�@�v�d�z߈� ��x�4�������� �h�D�.�2� �$[�'G�[�^�B���B��CH� ^�� ��u�����������p�h�M�_�q�����T�����^�^��Y�m�2��
  ����#5GYk }������h*��� ��>�x}���$MSKCF�MAP  ��?� �����m�N"ONREL7  6�9_��"EXCFENB�k
7]�FNC��}JOGOVLKIMkduyd"WKEYk�"WRUN��"SFSPDTYU�x�v_SIGNk>}T1MOT�z�"_CE_GRoP 1n��9\���/���/�/4��/ ?�/2?�/'?h??�? C?�?�?y?�?�?�?O �?@ORO	OvO-OoO�O cO�O�O�O_�O*_<_�#_`_-�"TCOM_CFG 1o/����_�_�_
|Q_/ARC_�6��UAP_CPL�_��NOCHECK� ?/  5�;h9oKo]ooo�o�o �o�o�o�o�o�o#�5GTNO_WA�IT_LF'5y"NMT�Qp/���qo_ERR�!2q/_�� R_����"�:�L�dT_�MO�sr�}, �C�P_��_�PAR�AM�rs/�������MW��� =�e�345678901.�@�R�)�q��� _�����˟����ݛLW�3�E�؏i�c�UM_RSPAC�E,�������$ODRDSP�SI&��OFFSET_C�ARToݨDIS��ݢPEN_FI�LE�I!�Q�v�PO�PTION_IO����PWORK kt�'� T� |�C�����6���Z����	 �m���C�
����RG_DSBL'  ��v����ޡRIENTTO�j�C���8=�#�?�UT_SIM_DJ�6	���VàLCT u��}�����Q��W�_P�EXE���RAT����� ���UP� ve������`�����*�8��$���2�#h)deX)�dh�O�X dY�ߑߣߵ����� �����!�3�E�W�i� {������������2n��)�;�M�_�q� ����������<��� ��+=Oas@���X��� O���1m(���(��.�g��"0 �дu�  @D7�  �?���?р��D4  �EzZ3;�	�l	 0DӀS@SM� �i��i �H)!H�,�H8�H�m�G�	{Gǎ8��6�MV���� �C�)����)����Ճ�*�  �p  �z > �  ���/$"�,��B,�Btr�«���O¼�/���/��"�# �,0 �}� �  � �߽pj   ���&X�?MU	'�� � 12I�� �  ���-=���U?g;/�@}?�0~.ѱ�?�;Ѳ���H[N ��?A'M�D�> C%)�f)�" B& ��"O4B+�:�Q��@D1�oo�$�����JWAD0�J@�A: �1�E&?�O��O#__G_2]��� �t O�� ru �4� ��R�U���' :�%S�р�? �?�ff��@[�_�_V_{�o~��118р"o0j>�P�Q6YPрZo�WrAdS�%�>Lw0�#��<	�I<g��<5�<2��<D��<�׍�l��_�ѳMb�@?offf?�0?&p�:T@T�q?��`?Uȩ?X�-q�iyBq5Y a��gI�_� �����!��E� W�B�{���d�����Տ�LnpΏ/�ʈG�@ G��U�ȏy� d�������ӟ����� ��yB=� ��?p�� �/򏸯�߯R��� '�9��oN�`�����~�P����ۿƿ�B�� �D�e�ֿ;�ҿ_�J�?��h�oϨϓ�J���D4��b!�_@ ���� ߧ��Ŀ�����%�@I�)�M`�B@��@`��9@y��?��h	� �@�3��[N��N�N��E��<�/�Y�kЖ>��ڟ��A�p�C��F@�S���pX������@��t��%�h���߉!G��G�knF&�F׿�pE,8{�� �F�ZG����F�nE��DE,ڏ������G��F7���F��ED��Mf��b�M��q�� ����������(�� 8�^�I���m������� ��������$H3 lW�{���� ��2VAS �w������ /.//R/=/v/a/�/ �/�/�/�/�/�/?? <?'?`?K?p?�?�?�? �?�?�?O�?&OO#O \OGO�OkO�O�O�O�N=(]�3�ji�O�a���	U�E3Ա�x�O_�a4 ��%_<7_�a�P�Q_c_�ERjb}_�_1w?������]�Y��_�_o�_1ol��P�bPcn~���o�O@�o{_�o�oY�`��o �o,/;M#�f 0o�����Y�e@t�~�i#�1�C�yM� _�����������{bS� Ԏ��	�?�-�c�Mj�2���$�VG�Dz}�B����B��CH�}�9�֟��� ��0�B���wl�@~�������Ư�T�E��\��qQ��U
 ί�0�B� T�f�x���������ҿ����χ��� ���]{x}��$P�ARAM_MEN�U ?Յ��  �DEFPULSE��	WAITT�MOUTl�RC�V� SHE�LL_WRK.$�CUR_STYLvj���OPT��N��PTB����C��R_DECSNw� Te'�!�3�E�n�i�{� �߶߱������������F�A�USE_P�ROG %P�%�B��V�CCR���UeXÚ�_HOST7 !P�!����Tt`����������4���_TIME��� �T�  A�GDEBUG��P�V��GINP_FLM3SK]���TR����WPGA�� |�[����CH����TYPEM�Y�A�;�Q zu������ 
)RM_q �������/ */%/7/I/r/m//�/��/�/�/�/?��WO�RD ?	��	�RS��CPNeS�E��>2JO��ξBTE���TR?ACECTL�PՅ�Z� a`;/ <a`{`�>�q6DT QxՅ��0�0D�����0��2��2U�4�4	�4
�4U�4�4�4���Sc{a4@��:B��*O<ONO`HlE�0wB�0�B�?��?�?
OM�O�BkL_&_8_J_tO�Kl_ �K�_�_�_�_�_�_�_ 
oo.o@oRodovo�o ZO�o�o�o�o�o�o *<N`r���0����q�s���B��B��B��A �&��d�v����� �O�O�O�O�O�OЏ� ���"O�������� ��ƏH��1�] �2�D� V�h�z�������¯ԯ ���
��.�@�R�d� v���������п��� ��*�<�N�`�rτ� �ϨϺ��������� &�8�J�\�n߀ߒߤ� �����������"�4� F�X�j�|������ ��������0�B�T� f�x������������� ��,>�bt ������� (:L^p�� ����� //$/ 6/H/Z/l/~/�/�/�/ �/�/�/�/? ?2?D? V?h?z?�?�?�?�?�? �?�?
OO.O@OROdO vO�O�O�O�O�O�O�O __*_<_N_`_r_�_ �_�_�_�_�_�_oo &o8oJo\ono�oV�o �o�o�o�o�o"4 FXj|���� �����0�B�T� f�x���������ҏ� ����,�>�P�b�t� ��������Ο���� �(�:�L�^�p����� ����ʯܯ� ��$� 6�H�Z�l�~������� ƿؿ���� �2�D� V�h�zόϞϰ�������$PGTRACELEN  ���  ��������_UP �y�����������_C�FG z��������<��� �<�Z�l�<�$�DEFSPD {/���a�����IN~'�TRL |/����8Lԃ�IPE�_CONFI+�}>���<�]x�LID(�~/���GRP 1���������@��
=�[���A�?C�C
�XC)��B��r������dL�z�������� 	 �r�N��Ҩ�� ´����B������������A���> �6>7�D_�������� ='�=)���������	 B-��Q�M���  Dz����
��&L7p [�������/�6/!/Z/��
�V7.10bet�a1<�� B�=q�"`ff@���">����!=���͏!A>ff޷!@�ff�"�\�)�"D��?� � �!@�!� �!Ap�#W��h/??*?<?FK;�w����O/ �?K/�?�?�?�?O�? O>O)ObOMO�OqO�O �O�O�O�O_�O(__ L_7_p_[_m_�_�_�_ ��_ o�_$oo!oZo Eo~oio�o�o�o�o�o �o�o DQy{/�#F@ {yw}�y{ ջy�-������ /�Z?l?~?w���t��� ��я��������� O�:�s�^��������� ߟ�ܟ� �9�$�]� H���l�~����_ۯ� �����5� �2�k�V� ��z�����׿¿��� ��1�\n�j�|϶ �������	�4�F� X�j�c�χߙ߄߽� ���������)��&� _�J��n������ �����%��I�4�m� X�����ί�������� ��!E0B{f ������ H�Zό�Vh�ϴϊ ����� �2�D�V� O/�s/^/�/�/�/�/ �/�/�/? ?9?$?6? o?Z?�?~?�?�?�?�? �?O�?5O OYODO}O �O���O�OtO�O�O_ �O1__U_@_R_�_v_ �_�_�_�_�_"4F xBo|����o� �o�o//0/B/;�_ _J�n���� ���%��I�4�F� �j�����Ǐ���֏ �!��E�0�i��O^� ��N�ß՟������ �A�,�e�P�b����� �����o o2oTo.� hozo�o�����o��Ϳ �o
گ'�֯K�6� o�Zϓ�~Ϸ��ϴ��� �����5� �Y�D�V� ��z߳ߞ��������� �1��Uy��:� ���������	���-� �Q�<�u�`�r����� ������T�f� x�n�������� ����7"[F j������ �!//E/0/i/T/f/ �/�/�/�/�/�/?�/ /?A?l�e?w?&?�?�? �?�?�?�?�?OO=O (OaOLO�OpO�O�O�� ��*�O_@RdZ_�l_��$PLID�_KNOW_M � ����A�TSV �v��P�[?�_�_o�O&oo�#o\o�B��SM_G�RP 1��Z� d�I`�oo�$Cf�d����D��TPbj�oLk �f�o"~�U�o> n2T�~��� ��7�4���p�D� ��R���ʏ�������� ��6�
�T��*�����V�QMR�c��mT�EGQK? GR��(� #���[��/�A�S��� ���������$���� W��+�=�O������� ����� ���S�����ST�a1 1�j�����P0� @����E�ϲ��� ������M�0�B�T� fߧߊߜ���������@��7��,�m��2��9���A�<��z�A3�������4���������5)�;�M�_���6x���������A7����������8�(:L��MAD � ���� ��P�ARNUM  ��Ko���SCH
�
 �
��S+UPD��xaq|{��_CMP_�`�� <Pz '�U�E�R_CHK��a��Z���RS���_�Q_MO� �%�_��_RES_G����� ��v/ {/�/�/�/�/�/�/�/ *??N?A?r?e?w?J'��W,g/�?L%��? �?�?N#(��?OON# w�4OSOXON#��sO�O �ON# �O�O�ON#d ��O__N"V 1�x�Uua�@cX��P}p�P$@cW،P}��P@@cV��P��"THR_IN�R���pbA%d�VM�ASS�_ Z�WM�N�_�SMON_QUEUE ��eT��`Ȩ`�N��U�N�V�2`ENqD4a6/NiEXE]o�NeWBE\`>o/cO�PTIO;g?+2`P�ROGRAM %j%1`O_�0b?TASK_I��nOCFG �ox�9pDATAɓ]�B{@ev2w� �����z��+� =�O��s���������^nzINFOɓ��}�!dr��!�3�E�W� i�{�������ß՟� ����/�A�S�e�w�4҇ބ��| �98q~�DIT �B|ׯj~WERFL~h�wS~�RGADJ {�ƪA�  ,��?E�8��Q�IOR�ITY�W���M�PDSP�a�j�U��WvT�OG��_�TG���Rj��TO�E�P1�ƫ (/!AF�PE5 �~��!tcp��>%�!ud�?�!icm<�Q_���XY_<q�Ƭ=�Oq)� *������Op��������� ���<�#�5�r�Yߖ� }ߺ��߳������&�=*�PORT�a��OpA%�_C?ARTREP~`Ʈ>��SKSTA�X!*�SSAV`�ƪ	�2500H80A9u�T毙䕣�ƫ�����`X#�x$�6�m�URGEU`�B��A)WFP�DO�V�2�W�q�?Q��WRUP_DEL�AY �Ưe�RO_HOT�hwR%z�����R_NORM�AL�n��6SE�MI:y�QS�KIP���X%�x 	����� ���X%-;% [mE���� ���!//E/W/i/ //y/�/�/�/�/�/�/ ?�/?A?S?e?+?�? w?�?�?�?�?�?O�?�+O=OOO1U�$RB�TIF��NaRCV�TM�����m@DkCR����A�<]h�BQ���A�T�=���@�>�)�|���������c��_�@	��I<g�<#��
<2��<D��<��
+__{_ �_)`���_�_�_�_�_  oo$o6oHoZolo~o i_�o�o�o�o�o�o�o  DV�_z�� �����
��.� @�R�=v�a������� ����׏�*�mN� `�r���������̟ޟ �����8�J�5�n� Y���}���ȯ����� A�"�4�F�X�j�|��� ����Ŀֿ�ӯ��� 0�B�-�f�Qϊ�m�� ���������,�>� P�b�t߆ߘߪ߼ߧ� �������(�:�%�^� A����ϸ�������  ��$�6�H�Z�l�~� ��{������������  2Vh��� �����
. @R=O�s�� ���/�*/</ `/r/�/�/�/�/�/�/��/??&?28�AGN_ATC 1��K� AT&�FV0E02;�ATDP/6/9�/2/9p8AT�A2>,AT�%G1%B960�k9+++�?,�1H�?,�AIO_TYPE  E�C/4?REFP�OS1 1� KO x�O[H/ O/�O�MNO`O�O�O �O_�OC_�Og__d_��_+K2 1� K LON_�_o�_*o�_5A3 1��_�_�_ o�o�o�o@oS4 1�Woio{o�o3W>�oS5 1��o�o�J���jS6 1�����]��H����S7 1� �(�:�t��ݏ���S8 1�����Ϗ�	���r���)�SMA�SK 1� O  q
���ɗXNO�?��1.�8�1AMO�TE  �.DN�_?CFG �U����5�0BPL_RAN�GQ�K!Y�POWE/R �Q5 a��SM_DRYPR/G %�%R����ȥTART �����UME_PR�Oׯ�d�.D_EX�EC_ENB  y�5]�GSPD=�p���Y3��TDB��洺RMÿ��MT_�ѐT��S�D0OB�OT_NAME ��S�;9OB�_ORD_NUM� ?��A/H80�0I$�_	��s	�\������ ��en��	@�}�D|���D0PC_TIME�OUT�� xD0S�232n�1�Q;� LTEAC�H PENDAN��j�5��=Q�x0�Mainten�ance Con�sK"-��"+�t4�KCL/C�}��6��|� No Use�=[߹�F���NPO�ќ�5��_���CH�_L@��U���	�J��MAVAI�L`���+��]�I�S�PACE1 2�=L ���وp��扢J@����8�?��� �� �V�w�N��������� ������4�&G
 l�}d	Q5U1����� ����`4&G
@l}d�#��2��������2 A/b/%/w/�//�/�3����	/�/-/ O/^??B?�?�?�?�?�4�/�/??&?�? J?l?{O�O_O�O�O�O�O�5�?OO1OCO �OgO�O�_�_|_�_�_�_o�6_*_<_N_ `_o�_�_�o�o�o�o�o!�75oGoYo ko}o+�o�o��� �)��>��8Rd v��H������ӏ%�F�-�[��G ;�� R�;�
�� ����ԟ ���
��.�@�����c���p���8�¯=�d ؠ��ϟ���!�3�E� W�i�_�q������x� �կ��'�9�K�]� oρ�w��ϛ���Ͽѿ ����5�G�Y�k�}� �ߡߗ��߻������w `S� @���8堯F�"�*ل�� ���߇����� �,����V�h�2�<� N������������� .L4v�R\ n�����
f�7��_MODE  y��MS ���&����Ïb���*	�&/�$CW�ORK_AD]���x�!R  ��t +/^ _I�NTVAL]����hR_OPTIO�N�& h�$�SCAN_TIM�\.�h�!R ��(�30(�L�8������! ��3��1�/@>�.?���S22��411d�8�1�1"3��@���?�?�?h���IP���@���JO\OnOE@D���O�O�O�O �O�O__(_:_L_O���4X_�_�_�8�1��;��o�� 1��pc]�?t��Di�1>��  � lS2�� 15 17oIo[omoo �o�o�o�o�o�o�o !3EWi{�� ��wc���	�� -�?�Q�c�u������� ��Ϗ����)�;� M�_���`[����ğ ֟�����0�B�T� f�x���������ү������$�7�  0 ��� om�������� ǿٿ����!�3�E� W�i�{ύϟϱ����� ��v���/�A�S�e� w߉ߛ߭߿������� ��+�=�O�a�s�� ����ߖ����� �� $�6�H�Z�l�~����� ���������� 20DVP�\�  �A� ������ %7I[m��������/ �/C(/N/`/r/�/ �/�/�/�/�/�/?Fa;/?B?F�x1� ;?w=	12345678{_��l�@�P�?�?�?�?�?O9/2ODOVOhOzO�O �O�O�O�O�O-/
__ ._@_R_d_v_�_�_�_ �_�_�O�_oo*o<o No`oro�o�o�o�o�_ �o�o&8J\ n���o���� ��"�4�F�X�j�|� �����ď֏���� �0�B�T�f������� ����ҟ�����,� >�m�b�t����������ί����(��6 yI�[�@�`����������Cz  Bp�*   ���2�54F��$SCR_�GRP 1�(��e@(�l���0@ >`1 [1s�	  )�3�C�<�t�vrY��8P�}�kϤ���-�95C����-u���ȡ���LR� Mate 20o0iC �190�1�Շ0LR2C ��3�=OÆ�D�
f؜1u�2�U7��`1���v��@�u���	�t���������$�^0�2���_2T�g� �ϊ��o�F�D�f?��s�����￶ht ,�Z��sЬN�B��˰�P�N�g�N�Aܰv�  @DЎ�N�9@����  ?� ���J�H˰��y�N�F@ F�`������ A,Qwb� ��n�N�������B��_ J�n����� /�%//I/��E+:3 ��6?|?�5��
�/�/��#��@=��"��/pǢ� 3B�07��590@7���E�L_DEFAUL�T  I����� ^1MI�POWERFL � V�v5]2�0WF�DOk6 v5 �E�RVENT 1����O�t3C�L�!DUM_EI�P?�8�j!AF_INEj0O�$O!FT�?=NOraO!Q�O �PO��O!RPC_M'AIN�O�H��O�ON�CVIS�O�I��O�E_!TP8PPU�<_�9d4_�_!
P�MON_PROX	Y�_�6e�_�_XR�_��=f�_)o!RD�M_SRV*o�9gouo!RR8�o�4Yhdo�o!
�@M�_��<i�o!RL�SYNC4y8|�oY!ROS�?�|�4H�tO�8c �����;��_� &���J���n������ ��ȏڏ7�I��m�4��X����7ICE_�KL ?%�; �(%SVCPRG1�����!��3*�/��4R�W��5z���6�����7ʯϯ�C��5�9��oG���� o������D���� l��񑔯�񑼯7� ��_������4� ���]��������� ��'��տO����w� �%ϟ��M����u� ���������?�A� �Ͽ�ђ�؟ꐊ��� ɱ��������?�*� c�N������������� ����);_J �n����� �%I4mX� |�����/� 3//W/i/T/�/x/�/ �/�/�/�/�/?/??�S?Ś_DEV ��9�MC:�[8�im4OU�T_Rf1~6i8RE�C 1���f0�0� f0 	 �f0�2  
f0��4�1���3OMK��1�4=A%O^OAA��
� �Z�6 s;B�3AAqE=�=AP���2WG�1f0)f0�{f0U�Of2B0�O����/Q0�OP_�5��@��@r�H}�;@�  x�0�}@U@��O Rf0�f4�1af0�V_��2X0��@�f0?b�@�~_�__��2\��0��0��0�@�����_ f0�Tf0�1=f0[f0�o��2T0��@�f0*b�@u*oco�_�ÆL�H�0�0��R �  �RobmU�f0zf0�o�2�QU��@�f06�@z�o�vo~K�L=A�1(�f0tf0�f0�_c�hf4e�=�ZZ f0Uk0��0Cf0f01q��"~N�LiIP�1�2�f2Pf0>jIT��zDf0f0o.��g���φL"f0i��0bf0��0��0TV�b�f0f0/f0M|~ 0��E0��@�f0$�@Y�^�p���ՆL*�A�0=њQpɀ��b�Jʈ�f0_^�f2C0%��@��A0�����&��2\�AM��FUp��A��p�<~��O��Ӧ�$2�k�ҟK�2\&f0}��0+�0Wf0�Z��bU�f0f0R~�[��J�F��@ݒq0"ޯ �*�a@��Z�H� ~�l�������ؿ��� ���2� �V�D�zό� nϰϞ����������� .��>�d�R߈�v߬� �����������*�� :�`�N��f�x��� �������&�8��\� J�l�n����������� ����4"XFh �p����� �0B$fT�x�����5V 1a��<���0��O��2k0��0��>a?_TYPE�?k2�HELL_CFG� �z:f2/ qHL�/<7RSա �/�/�/"??F?1?j? U?�?y?�?�?�?�?�?`O�?0OBOQK��p�!%QOO�O%��x��q�qQ��M�q�pވ"(hAQ�d�O�O�&H�K 1��+  �OE_@_R_d_�_�_�_ �_�_�_�_�_oo*o�<oeo`oro�oa&�#OMM ��/�o�"FTOV_ENM��t"!}*OW_RE�G_UI�oe"IMWAIT�b���G${�OUTv$&yT�IMu��`V�AL5's_UNI�T�c�v})MON_�ALIAS ?e~�i ( he! � ��$�6�%��c� u�����D���Ϗ�� ���)�;�M�_�q�� ������˟ݟ���� %�7��H�m������ N�ǯٯ������3� E�W�i�{�&�����ÿ տ習���/�A�� e�wωϛϭ�X����� ������=�O�a�s� ��0ߩ߻����ߊ��� �'�9�K���o��� ���b��������#� ��G�Y�k�}���:��� ��������1C U y����l ��	-�Qc u�2����� �/)/;/M/_/
/�/ �/�/�/�/v/�/?? %?7?�/[?m??�?<? �?�?�?�?�?�?!O3O EOWOiOO�O�O�O�O �O�O�O__/_�O@_ e_w_�_�_F_�_�_�_ �_o�_+o=oOoaoso o�o�o�o�o�o�o '9�o]o�� �P������s��$SMON_D�EFPRO ����:�� *SYS�TEM*  �l��*�RECAL�L ?}:� (� �}7copy� virt:\o�utput\ca�lprxy.pc� md: ove�r =>1724�25216:46�795 432 ?291652�͏Lߏ�s}6z���z�������B�T��y�\toest_��ls�ਏ:�˟ݟ��!er�srch 0x1_60002�� �� ��?�Q�c�v�����,� ��ϯ��������M�_�򏄪z��$�6� ǿٿ���&�����?� Q�c�v�����,Ͻ��� �����Ϫ���M�_� rτϖ�(�:������� �ߦ߸�I�[�n߀� ��$�6���������� ���E�W�j�|�� � 2����������	��ASe}4z������%�/��� };z� �tp~� -��GYl�	��#�1��g?�	� %���L/^/q���@��3/�/�/iA� ��	/6�/,<?N?`?�stpdisc� 0=>lapt�op-3jv24�8ms:16104 ?,?�?�?�?t�tpconn 0 �?�?�?�?JO\O�o
xyzrate 61 OO)O�fO�O�O��zG�?30348 �O�O?_Q_ c_v?
__,_�_�_�_ �?�_�_�_;oMo_o�
�frs:orde�rfil.dat���tmpback�\�_S6o�o�ol2>�b:*.*�o�o@P�o>Pbuxzd:\�pS1��g7zua��X �C�U��z/�� ��3P0144:6949731�ԏg�y��z������B� T��y��/�����ҟ ��/	?�N!�<�N�`� �����1�¯ԯg� �~�*���L�^�qo �o\6�ǿٿ�o�o���"��E�W�f��$�SNPX_ASG 1�������� P �0 '%R[1]@1.1f���?��%���Ͽ�  �����6��@�l�O� ��s߅��ߩ�������  ���V�9�`��o� ������������� @�#�5�v�Y������� ��������< `CU�y��� ���&	0\? �cu����� /�/F/)/P/|/_/ �/�/�/�/�/�/?�/ 0??%?f?I?p?�?? �?�?�?�?�? O,OO PO3OEO�OiO�O�O�O �O�O�O_�O _L_/_ p_S_e_�_�_�_�_�_  o�_�_6oo@oloOo �oso�o�o�o�o�o�o  V9`�o �������� @�#�5�v�Y������� Џ��ŏ���<�� `�C�U���y���̟�� �ӟ�&�	�0�\�?� ��c�u��������ϯ ���F�)�P�|�_��x�PARAM ���� ��	���P���p�OFT_KB_?CFG  �����״PIN_SIM  ��̶�/��A�ϰx�RVQST_P_DSB�̲�}Ϻ���SR ��	�� &  E�ST_MV�����ԶTOP_ON_�ERR  ������PTN z	��A���RING_PRM��� ��VDT_?GRP 1�����  	з��b�t� �ߘߪ߼�������� +�(�:�L�^�p��� ��������� ��$� 6�H�Z�l�~������� �������� 2D V}z����� ��
C@Rd v������	/ //*/</N/`/r/�/ �/�/�/�/�/�/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4O [OXOjO|O�O�O�O�O �O�O�O!__0_B_T_ f_x_�_�_�_�_�_�_ �_oo,o>oPoboto �o�o�o�o�o�o�o (:Lsp�� ����� ��9��6�׳VPRG_CoOUNT��ќ��d�ENB/�_�M���鴖�_UPD �1�	�8  
 M�������-�(�:� L�u�p���������ʟ ܟ� ��$�M�H�Z� l���������ݯد� ��%� �2�D�m�h�z� ������¿Կ����
� �E�@�R�dύψϚ� ������������*� <�e�`�r߄߭ߨߺ��������\�YSDE�BUGn�Ӏ� �d���"�SP_PAS�Sn�B?4�LOoG �΅��� ���
�  ���� �
MC:\x`��a�_MPCf�΅����ҁ��� �ҁ��SAV �bi���� ����SV�TEM_T�IME 1�΋� (   ��	����T1SV�GUNSɀo�'������ASK_OPTIONn�΅�������BCCFGg �΋O� H�2!`;A�I�r ]o������ �8J5nY� }�����/� 4//X/C/|/g/�/�/ ��,�/�/ ??�/ �/H?3?l?W?�?��? ��0�?�?�?O�?&O OJO8OZO\OnO�O�O �O�O�O�O_�O _F_ 4_j_X_�_|_�_�_�_ �_�_o�X�  o2oPo boto�_�o�o�o�o�o �o�o:(^L �p����� � �$��H�6�X�~�l� ����Ə���؏���� �D�2�h�o������ ԟR�����.�� R�d�v�D��������� �Я����<�*�`� N���r�������޿̿ ��&��J�8�Z�\� nϤϒ���~������ "�4߲�X�F�hߎ�|� �����ߤ������� B�0�R�T�f����� ����������>�,� b�P���t��������� ����(��@Rp ������� $6ZH~l ������� / /D/2/h/V/x/�/�/ �/�/�/�/
?�/?? .?d?R?�?>�?�?�? �?�?r?OO(ONO<O rO�O�OdO�O�O�O�O _�O__&_\_J_�_ n_�_�_�_�_�_�_�_ "ooFo4ojoXozo|o �o�o�o�o�? 0 BT�oxf��� ������>�,� b�P�r�t��������� Ώ��(��8�^�L� ��p�����ʟ��ڟܟ �$��H��o`�r��� ����2�دƯ�����2��P��$TBC�SG_GRP 2���� � �P� 
 ?�  {���w��� ��տ��ѿ���/�A��T�[��b�d0� �p�?P�	 H;BHA�L�͌�@�B   C���϶˘���ϟ�D����AQ���x���A��T$��9��6ff��f�@2P�C�ώ�@�f߬��C��ߐ߮ߴޥ� ��%��%�D�W�"�4��j�|�������?�Y�����	�V3.00s�	�lr2c��	*�2�*�O�A� ��ѳ3e3P�d��� x�J�y�  �������T�JCFG Ė�l� o������������=K
%�Kq \������ ��7"[Fj �������!/ /E/0/i/T/f/�/�/ �/�/�/�/s���?? (?�/[?F?k?�?|?�? �?�?�?�?O!O3O�? WOBO{OfO�O�OP�<� �O��O�O�O0__T_ B_x_f_�_�_�_�_�_ �_�_oo>o,oNoPo bo�o�o�o�o�o�o �o:(^L�� ����h� ��$� �H�6�l�Z�|����� Ə��֏؏� ��D� V�h�z�4������� ҟԟ��
�@�.�d� R���v��������Я ���*��:�<�N��� r�����̿���޿ � &��>�P�b�ϒπ� �Ϥ϶��������4� F�X�j�(ߎ�|߲ߠ� ����������B�0� f�T��x������ �����,��P�>�t� b��������������� &(:p^� ���t����� 6$ZH~l�� �����/2/ / V/D/z/�/�/�/j/�/ �/�/�/?.??R?@? v?d?�?�?�?�?�?�? �?OO<O*O`ONOpO �O�O�O�O�O�O_�O __&_\_�t_�_�_ B_�_�_�_�_�_"oo Fo4ojo|o�o�o^o�o �o�o�o�o0B�o xf����� ����>�,�b�P� ��t���������Ώ� �(��L�:�\���p� ����ʟ��� ��_� *��_�l�Z���~��� ��į�د� �2�� �h�V���z���¿Կ 濠�
�����.�d� Rψ�vϬϚ��Ͼ��� ���*��N�<�r�`� �߄ߖ��ߺ������ �8�&�H�n�\��� >�����x������4� "�X�F�|�j������� ��������
T fx�D���� ��P>t b������� //:/(/^/L/n/p/ �/�/�/�/�/ ?�/$? 6?��N?`?r??�?�? �?�?�?�?�? OODO VOhOzO8O�O�O�O�O��O�N  PS� V$_R�$T�BJOP_GRP� 2��E�  ?�W�<RCS�J\��@'0WP�R@T�P� � ��T�T� �Q[R	 �B�L  �UCр �D*W[Q�_�_?f�ffe:lB} �P�ff@`�33D  $a �U3o>g�_�_po�l�Pޔe9<�bbY��?٪``$o�oU�A��gD�`$��co�Quz9�PӜAa�P@a�̇�C�Z`Ep�o]Ag6ffpu`aD/�U�h�͔r��~�a��RieAq�`�q��@9q�|�d&`%��΃c333D�\P8�7��?�`?L�pAp[QB�b�k�}� ��|z�� >�ffԁL���T�f��fo  ��Nw@�*�8�f��� r�,���П��ȟ��'� ���F�`�J�X������SC�Vء��	�V3.00�Solr2c�T*��TQ�� E����E�A E���E��3E��iNE�!hE��فEۑ�E��I�E��E����E�rF��F�F�M(F�5F�BFaOF�\F"f,��z  E�@ E��� E�� Eߙ  E������ E����� E�Ȇ�Ԏ�ᆰ�� F   F�� F$ Fj`� F�@ F�P� F�` 9�I_R9�o��赢L�_ ��V���LQ�8TESTPARS�XUP9S�HRk�ABLE K1�J[4�SVȢ+� �0�V�V�PV�WQV�	V�
V�QVȥ�QV�V�qV�뱅�RDI��TQ�϶���������f�On߀ۊߜ߮���$�ކ�Sl�RS 0ړ� ������������#� 5�G�Y�k�}������� ������/]k�o��*	 �%�7�I�����+��=�O؆�NUM [ �ETQ�P�P �밆�_CFG ����Q�@<PIMEBF_�TTq��RS~�;V�ER�<Q;R� 1�J[
 8$�RP� �@5  ������ //&/8/J/\/n/�/ �/�/�/�/�/#?�/?�Y?4?F?\?j?|?{_��h@R
<PMI__CHANG R} �3DBGLVQ`�IR;Q�0ETHERAD ?�E;@�S �?�?TO�6V�0ROUTe�!JZ!�D�OwLSNMASK0HRSAA255.�E��O��O8TOOLOFS�_DIq��5IO�RQCTRL !�s[���n]8]_�_ �_�_�_�_�_�_o"o 4oFo�
�_Tofo�og��PE_DETAI�H3ZPON_SV�OFF)_�cP_M�ON �"P2��iSTRTCHK� �J^mO�bVTCOMPAT�h�;C�d�`FPROG� %JZ%TP?REC T-=�m�%QPLAYr��j_�INST_M�@ 2�|�g�tUSe]�orLCK��{QUICKME�0)�oroSCREF�3Jtps��or�a�f��2w�_{���Zy�ISR_GRP �1�JY �� 6�����;�)�_�M��8���� Y�������͕��� ��/��S�A�w�e��� ����ѯ��������=�+�M�s�	12?345678�����f�X`�1�Ћ
 ��}ipnl/�۰gen.htm������0�B�X��Panel s/etupF�}<��`�Ϫϼ����� u� k��*�<�N�`�r��� ��ߺ��������� �ߝ�J�\�n���� �I�?������"�4� F���j���������� ����_�q�0BT fx����� ��>�bt�����3�~UA�LRM�pG ?J[
  �*/ !/R/E/v/i/�/�/�/ �/�/�/�/??<?��SEV  ��n6�ECFG ���m�6��A�1 �  Bȩt
  =?�s3E�?�?�?OO +O=OOOaOsO�O�Gz1ʂ��k SΟ�O�H7Isv?}{�`(% 0?"_p_I_4_m_X_ �_|_�_�_�_�_�_o0�_3o�L� �M�O�AoI_E�HIST� 1��i  �(k` ��(/�SOFTPART�/GENLINK�?current�=menupage,153,1}o��o&�o�o,166�or���7I[r2a���,�2�p'��~71�y���������q)C��ue�dit�bTEST�h����#�5�@�R�e,2�o���������<W��c48,2����,�>��,ϟُ�_MVp�������í�)a�a)o���%� 7�I�ȓޯs������� ��Ϳ\����'�9� K�ڿoρϓϥϷ��� X�j����#�5�G�Y� ��}ߏߡ߳�����f� ����1�C�U����� ����������Я	� �-�?�Q�c�u�x�� ������������) ;M_q ��� ����%7I [m���� ���!/3/E/W/i/ {/�//�/�/�/�/�/ ?��/?A?S?e?w?�? �?�/�?�?�?�?OO �?=OOOaOsO�O�O&O �O�O�O�O__'_�O K_]_o_�_�_�_4_�_ �_�_�_o#o�_GoYo ko}o�o�o�oBo�o�o �o1?�ogy �����o��	� �-�?��c�u����� ����L�^����)� ;�M�܏q��������� ˟Z����%�7�I� ؟��������ǯٯ h����!�3�E�W�Bz��$UI_PAN�EDATA 1��������  	�} � frh/cgt�p/wholed?ev.stmc����ӿ����)  ri��.�Ip��F�X�j� |ώϠ�ϲ��Ͻ��� ���0��T�;�xߊ� q߮ߕ��������Bv��� (�? #4�@�E� W�i�{�������6� ������/�A���e� w�^������������� ��+O6s�l�� ������� ��1C�g �������L 	///?/&/c/u/\/ �/�/�/�/�/�/�/? �/;?M?���?�?�? �?�?�?0?Ot%O7O IO[OmOO�O�?�O�O �O�O�O_�O3__W_ i_P_�_t_�_�_�_�_ Z?l?o/oAoSoeowo �_�o�o O�o�o�o +�oO6s�l �������'� 9� �]�D����_o�o ɏۏ����#�v�G� �ok�}�������ş,� ������C�U�<� y�`�������ӯ���� ޯ�-�����c�u��� ��������T��� )�;�M�_�q�ؿ��|� �Ϡ����������7� I�0�m�Tߑߣߊ��� :�L����!�3�E�W� ��{�� ϱ������� ���r�/��S�e�L� ��p������������ =$a����}�r�����)�*��Vhz ������� �.//R/9/v/�/o/ �/�/�/�/�/?��������$UI_PA�NELINK 1����  ��  ���}1234567890_?q?�?�?�? �?�4��]?�?�?OO 1OCO�?gOyO�O�O�O��OYIY0:�M���[0  SOFTPART/GENA1�?CONFIG=�SINGLE&P�RIM=mainedit �OI_[_�m_YJ_$_M=wi?ntpe,1@_�_ �_�_�]�_$o6oHoZo looo�o�o�o�o�o �o�o
2DVhz ������� �.�@�R�d�v��� ������Џ����M� 0,  9P E�=Por?S�5�co :�{�^�������͟ߟ ��'�9��]�o� R����O�O�����Z1 �/�%�7�I�[�m�`C �������Ϳ߿񿀿 �'�9�K�]�o��L�� �э͙�S�������� ���#ߒS;�M�_�q� �ߕߧ�6�������� �%��I�[�m��� ��2����������!� 3���W�i�{������� @�������/�� Sew����.� ��|�#G* k}`����� �/�1/C/֤�͡� ۯ}����/�/�/�/�/ ?�2?D?V?h?z?�? ?�?�?�?�?�?
OO �ϝϯ�dOvO�O�O�O �OE�O�O__*_<_ N_�Or_�_�_�_�_�_ [_�_oo&o8oJo�_ no�o�o�o�o�o�oio �o"4FX�o| �����e�� �0�B�T�f����/ ���������ُ��� >�P�3�t���i����� Ο��O/�s/(��/L� ^�p����������?ܯ � ��$�6�ůZ�l� ~�������#O5OGO� � �2�D�V�h���� �ϰ�������u�
�� .�@�R�d�v�ߚ߬� �������߃��*�<� N�`�r������� �������&�8�J�\� n�������������� ��m�"4ßXjM �q������ BT7x��� ���A��//,/ >/P/C�t/�/�/�/�/ �/�/o/??(?:?L? ^?Ϳ߿�?�?�?�? �? OO�?6OHOZOlO ~O�OO�O�O�O�O�O _�O2_D_V_h_z_�_ �_-_�_�_�_�_
oo �_@oRodovo�o�o)o �o�o�o�o*�o N`r���� �m��&�8��\� n�Q���u���ȏ��� ���"���?�?�{���$UI_POSTYPE  �5� 	k��{��_QUICKMEN  ���j�����RESTO�RE 1ו5�  � �/
�2�D�h�mc��� ����¯ԯw���
�� .�@��d�v������� W���˿ݿO��*�<� N�`�τϖϨϺ��� �ρ���&�8�J��� W�i�{��϶������� �ߡ�"�4�F�X�j�� ��������ߋ��� �y�+�T�f�x����� ?�����������, >Pbt���� ��(�L ^p���I���� //��SCRE�ܐ?�uw1sc-�u2M$U3M$4M$5M$6M$�7M$8M!��USE�R/ 4/F"T. O#k�sW#�$4�$5�$6ʶ$7�$8�!��ND�O_CFG ض��  ,� ��P�DATE �)��None �V��SEUFRA_ME  
��&�,1RTOL_AB�RT7?��N3ENB�X?I8GRP 1��!��Cz  A��3�1��?�?�?�?��?FO"OG:ېU�x81g;MSK  �{5�Ag;N41%�a��B%��O��VI�SCAND_MA�XyEI�c8�@FAIL_IMGy@�f���#�8�@IM�REGNUMyG
��KRSIZyC,����$,SONT�MOUW0{D�%��VU�#�c�� ��P�2FR:�\�O � �MC:\XS\LO�G�VB@4 !��O�_�Q�_o
�z? MCV�_�SoUD10fEX9k�
�f�wV�2ۜ�z�p(��=��͓o��j�o�o�o�o�o �o�o 2DVh�z��KPO64_r?S�0��n6�u�Q0LI Q�z�x�qV�� �|f@�w��w =	�xSZV�~w����wWAI���DSTAT ܄�;�@�_ď֏�$���EP12DWP�  ��P G�/����q�AP-��B_�JMPERR 1�ݜ�
  � 23�45678901 �������ʟ��ϟ� �$��H�;�l�_�q�x���LT@MLOW��8�P�@�P_TI_X�(�'�@MPHASOE  53���CSHIFTUB1=~k
 <���O b��A�g���w���ֿ ���������T�+� =ϊ�a�s��ϗϩ��� �����>��'�t�K��!��#ޛ:	VS�FT1�sV�@MN�� �5��4 �0���UA�  B8*���Ќ�0p����b�Ҫ��e@��ME*��{D�'���q��&%��!�M�$�~k���9@�$~�TDINGENDcXdHz�Ox@[O��aZ��S����.yE����G�� ��2����������RELE�y?w�^_�pVz�_ACTIV����H��0A �`�K��B#&��RD�p���
1YBOX ���-����2��D�190�.0.� 83���254���2�p�&��robot����   pxN g�pc�  �{�v�x���^$%ZABC�3�=,{�낆;-!/^/ E/W/i/{/�/�/�/�/ �/?�/6??/?l?!	ZAT����