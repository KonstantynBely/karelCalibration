��  ë�A��*SYST�EM*��V7.7�077 2/6�/2013 A�Q  �����ABSPOS_G�RP_T   � $PARA�M  �  �ALRM_�RECOV1   $ALMO�ENB��]ON�iI M_IF1� D $ENA�BLE k LA�ST_^  d�U�K}MAX�� $LDEBU�G@  
���A�PCOUPLED�1 $[PP_�PROCES0 �� �1��UR�EQ1 � �$SOFT; T_�ID�TOTAL7_EQ� $,�NO/PS_SP�I_INDE���$DX�SCRE�EN_NAME ��SIGN�j��&PK_�FI� 	$T�HKY�PANE�7  	$DU_MMY12� ��3�4�GRG_�STR1 � �$TIT�$I��1&�$��$�$5&6&7*&8&9'0''@�%!'�%5'1?'U1I'1S'1]'2h"�_S�ASBN_�CFG1  8� $CNV_J�NT_* �DAT�A_CMNT�!?$FLAGSL*�CHECK��A�T_CELLSE�TUP  P�� HOME_IO�� %:3MAC{ROF2REPRO8^�DRUNCD��i2SMp5H UTO�BACKU0 �� �	DEVI�C#TIh�$5DFD�ST�0�B 3$INTER�VAL�DISP�_UNIT��0_�DO�6ERR�9FgR_Fa�IN�GRES�!Y0Qy_�3t4C_WA�4��12HGX_D�#�	 d $CA�RD_EXIST��$FSSB_�TYPi� CHK�BD_SE�5AG�N G� $SLOT_NUMZ��APREV��|G �1_EDIT1_
 � h1G=�H0S?@f%$EyPY$OPc� �0LETE_�OKzBUS�P_CRyA$�4�FA^Z0LACIwY1�KR�@k �1COMM{ENy@$DGV�]QP� ��OF��BL*OU�B , $�1V1�AB0~ OL�UR�"2CAM_;1� x�f$AT�TR��@0ANN��@�IMG_HE�IGHyAcWID�TH�VTCYU��0F_ASPEC�yA$M@EXP�;$� Mf�CF�cD X $GIR� � S!1U`BfP�NFLIC`~d
U�IREs3��AOM>qWITCH}cX`�N.0S_d�SG0� � 
$WAR�NM'@f��@� L�I? �aNST� C�ORN��1FLT�R�eTRAT@0T��`  $AC�C�1"p '|�'rOcRIkP�C�kRTq0�_SF� 4 �CHuGI1 [ �Tz`u3IPpTYPVD�@*2 �P�`�� 1zB*HD�SJ�* ��q2�v3�v4��v5�v6�v7�v8��v9�CO�$ <� so�o�h�s1�P�O_MOR./ t 0Ev�sNG�8`TBA�  5c���A�����]@�!���ϋP�0Ѕ,*��h�`
P�@��2� �,p�J,p_!Rrrqo@+�J/r/�&J�JVq@�Cj��m��g��ustP_}0O�F� 2  @� RcO_���WaIT8C���NOM_�0�1�ەq3� ��cD Ԑ;����hP���mE!XpG�0� F�p%r
$TFx�JF��D3ԐTO�3&@U�=0�� �H,�24�T1��E�� �e��f��f��0�CPDBG;a� 6k@$�PPU�3��f):��A�A�X 1�dUN�$AI�3BUFuF����!� |�`��`PIV��Pr�Mq��M~�䠁�Fr�SIMQS��G��QE�ڿ�~��MC{� �$}1JB�`S�}1GDEC������ܴ�z� ě0CHN�S_EMP�r$Gg�=Ǎ@_��q3
p�1_FP󔞡TC h�@`�b��q0�c}�y�G�� V�AԂ�!!����JR!0ԂSEGF�RA.pv 7aR�T�_LIN�C��PV!F������Y����Q��)B����( '���f�e�S ���Q��.0�p�B��A����SIZC�ћԂz�T��g������QRSINF3��p�����?�������؉���Lpot��G�*�CRC�eFCCC�`+���T�h� �mh�SbA��h�*�f�D�:�D�d�c��C��PTA����w@�撀���EV���jF��_
��F��N&�G�� X�Y�����1i���! ��,��hRGNP��0qF���R}�qD���2}�LEWN� �Hc6���C�K��AA�>dCx :�L���ou2���A6N`CNo�$LGp��B�1 aP��s@�dWaA?@����~0R���dME`%`��d�_RAs3�dAZC���z�OFkqFC�RH`X`F�`p��}��,�ADI ;� 6b� ���`�p�`5cn�S�@1�7a&�AMP���PY8CU�IMwpU��iQU� $�P��C�CG1�������DBPX�WO����p$�SK��2(�DBT. TRL�1 ��Q0aTi� �P�DJ�4LAY_CAL�10R !'PL	3&@�0ED�Q5'ֱ5'̡����1!�W�PR� 
�1 0Δ1" �PA$��q$�� �LB�)#�/�#mp�0$�/��$C�!%�/�$ENEqr�&�/�#d �REp�"'H ��O)@"$LF3#$�#xB� W;����FO[ _D0m�RO(@���u��j���3�RIGGER�6P�A%S���ETUR�N�2RcMR_��T�U�`?�u0EWM����GN�P��zB�LA��E��$$EP#�CP� ��&@Dֱk�C5D�mpD�A�#�p4\1i�FGO_oAWAY�2MO��tfQg�CS_7(<�QIS � ���c�C���A����B�t�Cn��A"�F9W���DNTV@��BVkQ�����S˳W�s�U�J&�U�� ��SAsFE�ZV_SV6b�EXCLUl���N��ONLA��SY���Q�tOTBa��HI�_V/M�PPLY�_�a��VRFY_�#�q�Bd�_ �)0���_+�Ip� �TSG3� *�b݀�0 AM��� a*����0��Vi.b>%fANNUN� r�LdIDp�U�2~S @�`mijarj�f�P��堫@I�"+��c$FOb�׀OT@�w1 $DUM�MYֱ�d[!�d١��& �E, ` 8�HExs��b�S|B$�SUFFI��@ ��@�a5��g6�a�MSW�E- 8��KEYI����TMZ1^ӌqL�1�vIN��%�D�. D��HOST? !�rְ�t[ `�t٠�tYp�pEM>����$��SBL��UL��/ �|3�ίr�DT50�!0 ϴ $9��ESAMP�ԕF���������I�0��$SUBe�Q�� �C�:��G�SAV��r����G�C� ˇ�PnfP$�80E��YN_Bn�1 0��DIadb�@O���}$]��R_I�� �E�NC2_ST � 2
ԇ J���L�q~S�`;����!3�M�I��1:�p�4  AL�3�M��0�0K�4x'a��AVER�q8��}�M�DSP�v��PC�U���\�ެ�VALUŗHE4� ��M�IP@����OPP7  �THS ���6�S�F�	F􁳠dL�0�T���SC�Q�d:�ET�o�5zrFULL_DUY�da�0��O�w�h�OT���0�NOAUTO�!6��p$�\���cTl�
�C` �C����۱�L�� _7H *�L���n�b���$�0P�˴ ��ֲ��[!���a��Yq���dq��7��8��9R��0����1��1��U1��1Ⱥ1պ1�U1�1��2
�2�����2��2��2Ⱥ2�պ2�2�2��3J
�3��3����3��U3Ⱥ3պ3�3ﺕ3��4
�[���SE�"8 <��~��`�;I�����/��Q�FE�0�0� 9 ,���Q?hpz@^ ?(�А��ER@#��`!�A��� :�`$�TP�$VARqI�<��UP2�P3; �pq�TD��S�|�1`3�����r�B;AC�< T�pr���)��bP��@o�IFI)�@���U���P��QF�0��� =t ;'�Ԡ��P'�ST(&�� HR�&�r0E����	%�C��	���_Cr�N�r���B��p�h�FORC�EUP%bn�FLUS�`HN �E�h�^�RD_CMK@E(����IN_��&vP.g�REMM�F~Q��@���� 3
K	9N0�EFF���N@IN�A��OVM�l	OVAl	TRO�V���DT��mDTMX���m{@�
���? �*[ ��CL��_:p']@$�-	_
�;_T��X
���@AQD� ���}��}!V1� R�Q��LIMIT_Ƚa椀�M��CLmd}�RIV	�a���EAR��IO*P�CC�����B�Bg�C�M@��R �GgCLF�G!DYM(�/�aR#5TWDGЍ�| s% �SS& �s> P�a�!r1���wP_�!�(�!1R��E�3�!3�+5�&O�GRA���?w�i�kPW��ONT��EBUG)S&2*��p{@a�_E @� 2��QZ �T�ERMB5AK9OR�IG0BK5�U��SM_�Pr�G0C~K5���TA�9�DK5N �UP>B�E� -zAa��@.PY3.@A$S�EG�:f ELEUU�SE�@NFI,���2�1ޠp4�4B$sUF6P�$��FQ4@�wAG0T�Q�&�HSNST P�ATm�piBPTH	J�AߠE�p��2�P@؀	E)�؁��1R�@<�InaSHFT_��1|oA�H_SHOR �ܣ�6 �0$�7�@Dq�'�OVR#�na�@�I�@�U�b �QAGYLO=�z��I'"��oAj�!�j�ERV ��:Qh��J��OG @�B�0����U����R!P"�ASYM.�"��1#WJG�уES�A�YvR�U�T @���E)�ᥳEP!�WP!�W�OR @MB��GR�SMT�F�GR��3laPA.@��p|�q�uG � ����TOC�1�`P<�@ �$OP���P�pՓá ��O�񖌀RE�`RC�AOX�pтpBe�`RmE� u�h�A��e$PW�R�IM�ekRR_p�c4��qB H2�H���p_ADDR~��H_LENGqBPyqnq�q�R��S�I H��S���q0���u���u���u��SE��'�*�HS<��J $N�`���_OFF��rP{RM� Lr�TTP_�H�K; (^pOBJ?"ip���$��LE`C|!�ȠL � ��.��AB_~TS�s��S{`��*�LVN�K�R��eHIT��B-G��LO�qt�f�N�͂���`���`SS�{ ��HW��A�M��p`INCPU>�"VISIO������+��t,��t,��� _�IOLN��N̠��C�q$SLzQb��PUT_�$�`{�P �V�^��F_AS�"O��$L��I����A��U�0�@Af��`q�<PHY���ÓZ���sUO��#P `�� ����ڔ� �2�pP���`(�L��Y�B����UJ�Q�z�N�EWJOG-G��DISx�[�K-�f�#�R 
�WAV�ǢC�TR�CǢFLAG��"[�LG�dS �����Y�3LG_SIZo���������FD)�I�4�E� *��D0���c$��� 𖶦���K���D0��� SCH_��߅p��2��N��F�T����E�"~�������U�
�
�{`L�	�DAU/�EA�-��dE��;�GH�b;ᲐBO}O��Uh Aɒ���IT��y�[0ŖR;EC��SCR�𙃖ʑDIēS.@��RGO���˒����d��$����SU���W�Ĳ��Ľ�JGM$�MN�CH,�FNKEuY%�KM�PRGK��UFY�PY�FWDvY�HL��STPY��VY�@Y؀�Y�RS"��H1`uۺ�CT�� �R��� �$�U	�m�@��
R�ݠғ`�G=ن�@POd�ڻŦ�M��FOCUd�RG�EX��TUIK�I{�����	������I�M��@A�S�`��p�@������ANA����2�VAILl�C�L!�UDCS_H!I+4`�s_�Oe�
!"h�S���|�S����IGN4��F�J��9T�be�_BUj � �V !PT�$�*��rv�Ϥd�@�A
VrW !Pi�'��T�0�1?2?3?�_� X � �i�=a�5���Ņ�ID$� tbP5R�bOh �Ĭ\A�ST	�RF�Y�� �@�  W$E�C�y����8^�� Y L�؟ 0��@���`qFtǀ��FwҬ�_ Z i`����b����>0C��[ �p C�LDP	��UTRQ�LI{��T����F�LG�� 1�O�D�����LD���ORG������hW�>(�siT�r� 4\ A�#0��վ�Sy`	T�70#0' �$�!>�#RCLMC�$B/ T/�)Q��!=1I�p_dg] d�RQ73�$DSTB�p�  � 6��-8AX�R �/8I<EXCESH�bd�2Mp�1^��A2�Tt6��0_�p"6_A:&��;G?tY80K�d` \��GROU��t$M�B �LI9�CRE�QUIRDB�aLO�#KDEBUr� 1L
YM��agbʑ`@�4C�" 1ND��`�c`b���̨�CDC���IN'��C��Z`���H��N��a#�� ��EPST�� �c\rLOC�RITp��P�Ap�1� 1ODAQ��d MX��ON�cF� R�fV�	X��b�U����uu�FX0IG}G�� e �y @X�a��X�XR�Q%��Y	��X	��V<�0ғDATA$`�E�a��a�N��f t $MDEaI:�)Sf��^d�![g�H5P�@]ez��a_cANSW�a^d�a��^e�D�)ARz�� Xpg[ �0CU4�V�`��=URR2{�h �D2�`A��A�! ?d$CALI&0���GS�w2K�RINtb�t<�NTEg�(i�bCu��=RBqg�_N�qjPukr���$tht�2kuyDIV�&�DHi0jp+�l c$Vp�C�$M�$Z0R<!T 0R����b�emH ��$BELT˪ZA/CCEL���;�"�IRCO�݁m��yT���$PSi0
�L�0ڰW��Cp�8��T�9�PATH���.���3]��Pl1�_<�r��Ł�"S C�r��_MG��$�DD�9���$FW�`7`���.����DE�PPABN�e�ROTSPEEՂ@L� JN�@���(0��0$USE�_p�P&�ܦSYh>��p�! �QYN09A����OFFua��7MOU߁NGJ�܀sOL~�ٔINC�d�2Q��-2��� -2ENCSpa2U��,+4R�IN�I]�B����"n�VE��s^��23_UPօp�LOWL��[�` '���D>�2@Ep]�'��2C[pW�MOS����4MO��0�'P�ERCH  ��OV����蓼����� �$�8S+�� 2@����B��V�0^�O�L�0P��7O�U�UP"��������TRK��AYLOA�J��1���]�͵³3P� �RT1I�1	�� MO�O��-2�28 �`4�w�ٳ��?�pDUM2���S_BCKLSH_CW�P�ϐΦ� ���bn�"�y�Ñ���CLAL V��!���� ��CHK �SՐRTY����C�
�*!6a_�ä_UM�����C���SCL��W�LMT_J1_L< 0-օa:�E4�U�G�D�J�P�J�SPCd�ȑZ���3�PC �3�H_A@�2��C� cXT���CN_rN���.�S��%�V���:� ���W�9���C' �SH�r�*�*!9��9� p��^���9���P�A���_P��_ �"�Ŷ�!ճ����cJG����~�OG�׾,�TORQU��ON��޹*�B٢-�*�&L�_Wž�_�sj�P�sj��sj�Ir�I��%I�sFKP]�J�!��,c!�VC�0'4�2���1��{0��82��J�RK��+� DBOL_SM���"M�@�_DL�q�"GRV�q�j�sj�sKH_p��I���
COS��LN- ���� �p�	�p�	�����bFZ� ٦KMY��D�TH�eTH�ET0��NK23��s��s� CB�CB�sC&1n2�����s��SB�s��'GTS�1W�C.�2Q������$�'3$DU���8A!r���2P&��1Qb8V$NE�4�PI� ���"$%�v$�p�A��%p�'���LPH�5�"h��"S��3�3�3�"+3:2�pV��(V�(�p�,V�*V�;V;V";V0;V
>;VL9H�(�&�2�-�n�H;H;H";H�0;H>;HL9O�,OR�(O}I�.O�*O;UO;O";O0;O>;O2F�"�Y�T��'SPBALANgCE_T@SLE�H_�SPHq�hR��hR3PFULC�lX�R{W�R3Uz1i�
�UTO_����Tg1T2�Y�2N�� �`��Tq���Ps d���T�O�p!�L�INSEG���R�EVf��Q�DIF̨�zy1j_g�r1k���OBUa��t$yM�I`���SLCHW3AR>��AB��u?$MECH�TXˑ�a��AX˱Py�p�f�'�r�Pl 
�b�I��:�ROB�C�RW�-u��~�pMS�K_KP�tn P �P_��R��r_tn���18�c�a�_p`��y�_p�aIN:a�MTCOM_C��>�po  ݀g`~4�$NORES���r��`�rp 8fU�GRJ��eSD� �ABג$XYZ�_DA�!F�r�DE�BU:a�q���pq �_P$��COD��� 1����`���$BUFINDXra�Hp"�MORRs/r $�qU&��Ɛu��ӑy�^��bG�i�s � $SIMUL��8��>�<��F�OBJEjP���ADJUSψA'Y_I��8�D����s�Ԑ_FIב=s�TZ��c����`@b�"�(�b`p0G�D���FRIW�d�Tg�R�O%�A�Eb񊰓�O�PWO> Vpt0>>�SYSBU0[�$SOP��I�����yU��b`PRUN�rڕPArpDٖ�b��.1�_OUTΑ�a��t$�IMAGҊ�\pv PDaIM���1�IN[ �0�RGOVRDY�˒����P�/�a�� L_`�PB�}����RB�ʇ ��MkᜪEDTb��` �N�@M���~В�]�SLjPVpu� x $OVS�LfSDI��DEX���q�����o��	Vb��N�A��'���,�'�D�M~�Ҥ_SETK�Vpv� @U�^��ep�RI��j�
q�_�}������Gqdà*� w� H\q�`��ATU}S<�$TRCx 8T�X�ѳBTMڷıI��P�4}Ѱ���.Vpx D\pE���β�0Ehbϱ�����ϱEXEհ����)=��f�ym�]p԰U�P�L�$�`6�X�NN���������� w�PG�uzW�UBñ�e��ñ��J_MPWAI[�P�&��LO7��pFA`���$RCVFAIGL_Cwq�p��R9� �p�c��(�}�"�-�A�R_PL��DBTqB��,��pBWD �f�pUM*�"�IG�87��Qc�TNLW�"�"}�Ry�iӻ�E������Hp��DEFSP>` { L\p�`���_��Ճ��UNI����Ѐ�RD��Rb k_LA`Pͱ���pUq|-�#��q�O���XPc�N�PKET��
��Pq�Uq}� h�ARSIZAE5p��=��u�S̀�OR��FORMAT�Pg�COנq�<b�EM�d����UX8��,���PLIb�Uq�~  $�pPO_SWI�`���Hq�AXG�b�AL_ So���A�rB���C�rD��$E6L���C_lі� � � ����r��J30 �r��TWIA4Z�5Z�6�rMOM��f��s��4��pB��ADf���s����PU�NR ����s�������Rt��� A$PI �&E�kqE�p-~- �-�WC�0$���&�9q�gE��eS/PEEDL@G�� ���Ծ����)�9�����)��	)���SA�MWPx�0�1��MOVD�H$_S`Y%nHk%_��1�t�2�t@����c�v��8�H�PxIN����������(�+(+G�AMM<Vu!�$GGETE�U�ٓD5�z��
�PLIBRv����I�$HIu�_�L�ݰpB�&E�(A�.� �&LW�-�&�, �)	6�&1��f�`j���� $PDCK���ٓ_�����E���b7��a4���a9�� $I��R�`D�c�b~�Ե`LE�qkq���8�1��0�Gq��`Vp��P/aUR_SC�R��A�r��S_SAVE_D��8Ex�NO5�C��y�6�8@ {$E�.{I��G	{I�@ �J�KP�q��H� � ��x"Mao���s ����d��6W2U�C�qy��L�0Rt� �k�F��aE��3�W<�@[�jQWg@5r�U��R�R��Sc2jQML"��[CL�W��M)A�Tr� � $P9Y����$W`�fNG�O�`�b� b�b#�HЈ��a� (���c��X�O����Z�e��ހRt� p䠰p�3+zO�O�OаO�O�a5�_�r� |�E�8@��>vs�>v@��8@_�kwVvy�EހPu%��"rB�\�P�"tP���PM&�Q}U5 � 8*��QCOU�1 �QT�H#pHOL<�QH�YS��ESe�qU�E�p.BZ�O�� � q�P���%��UN\ְ�Q ��OE��p� P2�3��AÔ�ROG�����Q2(�O}�2�������INFO�q� �#�e����RȾ�OI� (�0SLEQ�с�рi�C�{�ID��L��`� OK0�r��!E� NU�!��AUTTA�COPYqu�?��`@EML�NI�M�X�C���� Y�RGADJʵq�i�X�Q��$Pഖ�`��W��P��`�0�������EX8�KYC0b�ѪObpr�q���$�_NA9!�������`��?� � Q����POR�A�B�S�RV0�)a�Y�DI��T_��{������P�������5��6��%7��8y���S8BL�=�m�MC_F�p��PL9A8An�ȰR ��9��Ѽ��$iB�����d� ,�0FL�-`L�C@YN�[�Mz��C?��PWRc���L��!�DELA4��8Y5�AD�a� �QSKIP�� �Q�4�OR`NeT�Q ��P_4� �ַ@lbYp�� ���������Ƞ��@ՠ��������9�1��J2R� L�� m4*�EXs TQ%� ����(Q����p������p���RDCf� )�`��X9�R�p������r��A$RGE7AR_� IOT�2�FLG��vi��M%P9C��B�UM_����?J2TH2N'��O 1�����G8 �T00 �����M�lѺ`I�8��REuFr1�q� l�h���ENAB{�(cTPE�0�1���i� m���^QB#��:��"��(����2�ҙ���ߠ������&�3�Қ�7�I�[�m���&�4�қ�����������
&�5�Ҝ1�C�U�g�(y���&�6�ҝ�����������&�7�Ҟ�+=Oas�&�8�ҟ�����^&�SMSK�q�|���a��E?A��MO[TEF����a@0��(Q�IOQ5�qIc(P��POW�0L�� �pZ�����#p%�L��U�"$DSB_SIGN�1�)Q%���Cl��S2�32��b�iDE?VICEUS�,R>'RPARIT��D!_OPBIT`QY�OWCONTR;��(Q��O'RCU� M~DSUXTASKT3�N�p[0�$TATUF`PU#�0L�����p_,PC9�$F�REEFROMS8p��%�GET�0�WUPD(�A�2V"�P� J��� !>)$USA^���x6���ERIO�LP@bpRY�5:"_>@� �P}1�!�6WRK�I[D���6��aF�RIENDmQ�P�$UFw���0TO�OLFMY�t$�LENGTH_VTl�FIR�`-C�R�SEN ;IUFINtR]��RGI�1�ӐAITI��4GX�ӱCI�FG2�7G1`��Ѐ3�B�GPR� A�O_~ +0!�1�REЀ�E3�e�T�C���Q�AV �G(8��"J���u1~!  ��J�8�%��%m���5�0G4�X T_0)�L|�T�3H6���8���%r4E3GU�W$�P�W�R�TD�����T��а��Q�Tm�=$V 2����1����91�8�02�;2
/k3�;3�:iva�9�=i�aa�^S�jR$)V��SBV�EV'�V�BK�����&c��p��F�"{�@�2q�P5S�E��$.rRC���o$AŠFwP!R��Gv]U�cS'�� p7��rD3I�� 0�@DqV`��p�d`���PE0�@��=�
B5S!/� ��aRg�����R�6�N AX�!$�A�0L(A���r/THIC�1Y���h�t1TFEI��q�u�IF_CH�3�qI0�G�a�pG1bxf�з�m���S@��_J�F��PR�ֱ�S���Ԁ�d �$�SР�Z�GROU��̃TOT�t̃D;SP�JOG���#&��_P��"O������j��&KEP(�I�R����@M�R@�A	P�Qn�E^�`�!�[��SYS6��"[�PGu�BRK�B �.��pIq�p��M���΂��`AD�!̃9�BS�OC׆�NӕDU�MMY14�p@S}V�PDE_OP�#�SFSPD_OVR=���C����OR�CNm0�F�.����OV��SFR��pU���Fn��!#�p�C��A�"LCH�����РOV�s0��Wb�@M��ĥ:�RO�#�ߑ�_�p�� @�@�u@VER�ps0O�FSu@CV? �2WD6���2�ߑj2Y����TR�!���E_�FDOY�MB_CiM�D�B�BL�b>�f��attV"Q�240�/p��N�Gg�z�AM�x�Z�0���¿_M�~��"7����8$C�A�7�D����HcBK81��IO�5q���QPPAʀ=�"�M�5�͵���DVC_DBxC~� � 3"�Т�!��1�����3����pН�*���U�3��CAB ��2VӆPѣIP��c��O��UX�SUB'CPU�r	�S�P  P���90^SQ׹c��."~��$HW_C�А���S��cA�A�pl_$UNIT��l��ATTRI"���	��CYCL��NEC�A��J�FLTR_2_FI_�G(��9&��1LP�?�>�_S�CT�CF_��F_��6��FS8!����CHA�1�wᇲ�"v�RSD�4"�����q�_T��PROX��>�� EMy_ܠr��8d��a d���a��DIb0!�RAOILAC��9RM��CLOÐ C��Q*q���3q���PR��S�Q�pU�Cr�s 	��FUNC��@rRIN'PѸ0��u��!3RA��B ����8F�Ğ�WAR~���#BLQ����A��������DA����	����LD)0��Q1�q2��*q1TI2rQ�ǁ�p$xPRIA�1�"AFB�P�!�|ߠ�<`�R���MsOI��A�DF_&@؅�51��LM��FAށ@HRDY�4ORG6 H���A�0 �MULSE&@"�Q��a �G�	���m��$d$�1$1 ���0��߮� xm�EG0�̃�`ARހ���09�2o��z�A�XE�ROB�Wd�A��_�œSY������S�WRI�@s1��STR��� ��(�E�� !	%1��AB( �/&�a�ӰOT0v^�	$ߠARY�s�f"���S@	�FI���*�$LINK(���!�a_%#��%{q�"XYZp82�*�q�#OFF��R�"�"�(j Bဂj�4С��n�3FI��%7�q���j����_J���%��#�QO�P_>$H+5�3�PT�B\1�2C��i�D�U�&62�TURN��2r�5t!}��p��|7FL�`���m�0��%+*7�	� 1��. K�M�&8�2�Q�2rQ�#�ORQ ��G��-(�+p��z��� 3q�E"��T�GOV�@-A��M*�y�4 �E:�E@�FW�J� �G���D��o�*� � �A7�P��y��E�A�G`ZU:ZU�CG�ER�
��	6�E���B�TAFQ��)4����r'�AXУa2.q �c�W�c�W�c�W�p�Z �0�Z�0�Z%@�ZK@�Z ��Z
!�V� �Y� 
i � i� *i� :i� Ji � Zi� ji� zi�a�ioDEBU{�$v� u��;q��"F7O�n�CAB��6��CV�z� 
fr����u kњw�!�w�!�w�1�w �1�w%A�wKA�w��p\0��"3LAB"2�|EwЄ�҂�3 �z EERVEN�� � $q�_�NAǁ!_�PO�����` f�M�_M�RA��� d r T���ERR��L��~ TYi��RI�qV"0�S��TOQ�T)PL��T�Ѕ_��|��J � p�PqTl X���_V1�bP�Q���#�2�2+������/@��p��5��$W��V���VN�[�$�@�� �S����Q�	EHELL�_CFGN�� 5%�B_BASƴ�SRvp0�K� E�S��Jϐ1a�U%Α2�3�4�U5�6�7�8�RO���� � NL:�3ABn��АACKwv��)�o�pu0iႩ_PU2��COq��OU��P���ӕ�����T=P�_KAR�0&��REm�� P����QUE٩��@����CSTOPI_ALzs��� �T���� SEM[�w�k��Mw�y�TY��SO`��DI���Є�=��װ_TMK�MA'NRQζ� E���$KEYSWI�TCH��Ѱ��H=E��BEAT���EpLE����&�U���Fd�����SO_�HOM� O��REF�@PRi��R� ʞ�C@�O0�p EC�O���� _IOC�M�4M�k�5*8��'�O� D�!ۧH�U��;�M7��@��3FORCߣ�� �x����OMq �� @Etxk�U�#Po1B�O�o3�B�4x��NPXw_AS��� 0ݐ�ADD��(�$S�IZߡ$VAR\�TIPr�q�
G�A(ҷ��
�˨r�Ht�n�SV�XC�����FRIF�R��S0%�7�x���NFѲE�АO� x�PSI�ڂTEC*�%CSG%L=�T�"�0&�V�xD��>�STMT
�2o�P\�BW�@?��SHOWw��P�S�V� K�� ���A00�0�Q��KЀ��O���_���i���5���6��7��8��9��A����6������20��F��
 ���� U ����� ����0��P �J@��:�1G�1T�U1a�1n�1{�1��U2��2��2��2��U2��2�2�2 �U2-�2:�2G�2T�U2a�2n�2{�2��U3��3��3��3��U3��3�3�3 �U3-�3:�3G�3T�U3a�3n�3{�3��U454��4��4��U4��4�4�4 �U4-�4:�4G�4T�U4a�4n�4{�4��U555��5��5��U5��5�5�5 �U5-�5:�5G�5T�U5a�5n�5{�5��U656��6��6��U6��6�6�6 �U6-�6:�6G�6T�U6a�6n�6{�6��U757��7��7��U7��7�7�7 �U7-�7:�7G�7T�U7a�7n�7{�7��v��VP$�UPD���  �P����x�YSLO��� � ��հ���׆�QTAS�sTƠ��AcLU}U����CU�z�WFdQID_Lѳ��UHI�ZI�$F�ILE_Σ�T��$u�_VSA��� �h��+`E_BLC�K(�8bg�AhD_CPUQi��Qi���So�d_R1�ɢR ���
PW,�d� �aLA�S���c�a�dRUN5��a�d�a��d��5��a�d�a�d ��T�pACC����X -$&qLEN~�3t��&p�����Iѱ
�LOW_A�XI(�F1&q�T2�mwM��ɢ����Ip����Q�yTOR.��&p�{DW��s�LACE���&p�����_MAuйv�u�w�qGTCV�|��wTڱ �;�1�<ѷt��_��s���J����M��ӠJH����u���u2q�2��������s�pJKцVK~�か���3ՃJ0���JJv�JJ��AAL�P����4�5Xr;�N1B�N��	��tL�p_k����"p���� `5`GRO�U�PY�ӲB$�NF�LIC�ө�REQ�UIREv�EBU`V�"q���кp2����#pɖ!qxг�� �\��APPRՐC����p
!�EN�CsLOz�,�S_M �ȋ�A��u
!q��� 䣠MC�r;�XrN|�_MGц�C���,`��N��p��BRK���NOL������Rϰ_LI��է����	JޠѤP��p��p@���p;��pD��p6�K��8��v�"q���� ҒMr:q�l�Gqz�PATH v�������Rx�����m��pCNR�CA���է���IN%rUCh�pwQ�Cd�UM�!Yop�����QE:p��Gp�����PAYL�OAͧJ2LHPR'_ANqQ�L�`[��W�K�g���R_F2�LSHRё�LO�\�䱕����ACRL_�����޷C�rXrH�P"�$H��^�FLEX� q}J%u� :2 Dv�p4�K�GYq�pPbt|F1Kљխ׃@�������E� ���/�A�S�e�w� ����y���ф���蘏�����J�ÊT���X ����υ ��څ��[� ���
�� �)��;��D�V�h�z���J��� � �������Q�IPAT��ё��EL�4� �ؘJ���vߐJE��CTRޱ���TN��F�ɗH�AND_VBp��ѹP`�� $&�Fa2��K��ШRSWb�Y�j��� $$	M��}�R��E��Uw�H��sA�PH�����Q���A���P��A���Aɫ���j`��D*��DɫP��G�`1)CST��9!��9!N̨DY�`���|�Y� 鰋�KыǦ�J�ч�s�U�ХP��&�/��8�A�J�S�=��� ; �t�.R66N�/QOASYM����Ґ¹���Խ��ٿ_SH�����筈4��+�=�O�JV��h�p'CI����_VI��dHN�u@V_UN!I�ÉD���J҅�B �%�B�̦D�ųD�F�̀���������*Uc����X��H�`���XQEN� v�D	IɠS�OwT)YP���� ��I�1A �Q�äQ�`Bc�S`� � p�a.a� � ME����R'R�1TkPPT�0) ���Qz�~���0�Xa�	iT@� $�DUMMY1��o$PS_��RF���)$Pf�aLAƏ�YP�jb�S$GLB_T>mU�e��PpQ p���Q� �X	�ɗ`�ST���ߐSBR��M21�_V��8$SV_�ER��OÐ�c�cC)L�`�bA5�O�RTP�T O�P � D� �`OB���LO˰&uq9c�`r�0�SYSqADR��TP�PTCHb �� ,&����W7_NA���tz�ބS�TSR���l =��M�u `�ys�u~�s��s ����������� 0�)�T�"�5�~��� B����s�?�?�?DY��XSCRE)�pϚȐST[�s1}�P!��tY�r u_� Aq� T	� �`ob��a`�l��ҤԊ�g�c�O� ISb�c��TN�UE�TG� �ñjp^`Sq��RSM_iqmUU?NEXCEPlV֑XPS_�a����޳�p���޳R�COU�ҒS� 1�d�U�E�tҘR�b9�PR�OGM� FL�7$CU�`PO?Q��ִ�I_�PH�� �� 8џ�_HE�P�����PRY ?��`Ab_�?dGbOUS�� �� @�`v$BU�TT�RV`��CO�LUM��U3�SE�RVx��PANEԋ q��P@GE�U�<�F���q)$�HELPB�l2ETER��)_��m�A m���l���l�0l�0�l�0Q�INf��S�@N0�� ǧ1�����ޠ �)�L�Nkr� ��`T�_�B���$H�b T�EX�*��ja>�RELV��DIP>�P�j"�M�M3�?,iŠ0ðN�jae���U�SRVIEWq�S <�`�PU�P�NFI� ��FOC�UP��PRIa0�m@`(Q��TRIP>zqm�UNP�T�� f0��mUWA�RNlU��SRTO�L�u���3�O�3ORN3�RAU��6�TK�vw�VI�͑�U� $�V�PATH��V�CwACH�LOG����LIM�B���xv���HOST�r�!�R��R<�OB�OT�s��IM�� gdS)} 2����a����a��VCPU_A�VAILeb��EX
��!W1N��=�>f10?e1?e1$n�S��ۆP$BACKLAS��u�n���p��  fPC�3�?@$TOOL�t���_JMPd� �<���U$SS�C6>N�VSHIF ��S�P`V��tĐG�yR+�P�OSUR�=W�PRADI��P���_cb���|a�Q�zr|�LU�A$O�UTPUT_BMc�J�IM���2��=@�zr��TIL��SC	OL��C����ҭ� Һ�����������o�od5�?��Ȧ2 Ƣ���0�T���vy�DJU2��� �WAITU����n����%��NE>u�YB�O� �� c$UPvtfaSB�	wTPE/�NEC�р� �ؐ�`0�R�6�(�Q��� ش�SBL�TM[��q��9p����.p�OP��M�ASf�_DO�r
dATZpD�J����|Zp�DELAYng�JOذ��q�3� ���v0��vx��,d9pY_���	�7"\��Ѽ�rP? N�ZwABC�u� ���c"�ӛ�
N��$$�C��������!X`N�� � VIRqT���/� ABSf��u�1 �%�� < �!�/�/??0?B? T?f?x?�?�?�?�?�? �?�?OO,O>OPObO tO�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�o �o�o�o�o�o{� ���AXLMT�s���#  �tIN8&8qtPREO���+vupXuLARM�RECOV �)XrzujF ��%�!d ������7��I�[�m�~�, 
��/��vNG5� ��+	 =#�
�ڏ�� PPLIC�5�?�%upՁ�HandlingTool -�� 
V7.70�P/36 ��
�]�_SW2�D�F0<j�W� 43Y�J�|9�K�7DA7?�����
&�X�e	^-�None��J������ �T7��	�rP_�V�iu�6s��UTO�z"�,tTy.�HGA�PON� %��!.�U���D 1�y� t�x�����y.�K�oQ 1�{  Hp*������	����uq��"�" g�!��Hե�w��HTTHKY��"ٯ����u� ����󿽿Ͽ���� �)�;�M�_�qσϕ� �Ϲ���������%� 7�I�[�m�ߑ��ߵ� ���������!�3�E� W�i�{��������� ������/�A�S�e� w��������������� +=Oas� ������ '9K]o��� �����/#/5/ G/Y/k/}/�/�/�/�/ �/�/�/??1?C?U? g?y?�?�?�?�?�?�? �?	OO-O?OQOcOuO �O�O�O�O�O�O����TOĀ��DO_CLEAND���{S_NM  ɋ����_�_�_�_o��_D?SPDRYR�_��HI!��]@�_}o�o �o�o�o�o�o�op1CU��MAX � bTQNQS�sqXbTB��o�B���PLUGGpb�cWo��PRC4`B�P]klo^�r�O�r=o��SEGF;�K�+�6��_�_}��������ŏ�0�LAPZom�/��+�=�O� a�s���������͟ߟ|�6�TOTAL�v|�y6�USENUZ��g� HXL�NR��R�G_STRING� 13�
�kM,�S�
���_ITEM1��  n󝬯��Я��� ��*�<�N�`�r����������̿޿���I/O SIG�NAL��Tr�yout Mod�e��InpB�S�imulatedޕ�OutT��OVERRW` =� 100��In� cyclHŕ��Prog Abo�r^Õ�>�Sta�tus��	Hea�rtbeat��MH Faul����Aler���� �'�9�K�]�o߁ߓ��� ^S��^Q�� ������,�>�P�b� t��������������(�:���WOR 9���r���L������� ������*<N `r�������PO������ �9K]o��� �����/#/5/�G/Y/k/}/�/DEV� -�/�/�/? ?)?;?M?_?q?�?�? �?�?�?�?�?OO%O>7OPALT��^A ��8O�O�O�O�O�O�O �O__(_:_L_^_p_��_�_�_�_�_LOGRIxp��avO�_*o<o No`oro�o�o�o�o�o �o�o&8J\n�_*�R�ݦqo� �����(�:�L� ^�p���������ʏ܏�� ���PREG bNK��$�r������� ��̟ޟ���&�8� J�\�n���������Ϳ�$ARG_r�D ?	�������  �	$�	[��]���.��S�BN_CONFIOG ��L�K��F�CII_SA_VE  �k��b��TCELLSETUP ���%  OME_I�O��%MOV�_H��¿ȿREP��|��UTOBA�CK��V��FRA:\8�c �8���'`��q8�c�,�INIa@�8�^�,�MESSAGz������>��ODE_D��}��C���O� ��,�PA�US!��� ((O��J�\�F� |�jߠߎ��߲����� ����B�0�f�t�%�~*TSK  5�x�ϕ�/�UPDT����d����XSCRDCFG 1��;� �������&�8�J�\�n��� \�n���������� "��F��j|�����/e�2�GR�OUN����UP�_NAܰ��	�2��_ED��1
���
 �%-B?CKEDT-��}��p��Ѳ-(2�p8�/�/�8���g2���E/��/��/~/��ED3n/&/�/J/\.p�/"?�/�/ED4? �/?�/\.[?�?5?G?ED5�?n?#O�?\.p�?jO�?�?ED6ZO O�O6O\.�O_}O�OED7�O�Ok_�O\.pG_�_!_3_ED8�_�o�]-�_Vo�_�_ED9Fo�_�o"o�]-�o�oio{oCR oY_Vh�]1��{� LNO_DE�LGE_UN�USE	LAL_OUT V���WD_ABO�R���~�5�ITR�_RTN�ǀH�N'ONS)Ю������CAM_PARA�M 1����
 �8
SONY �XC-56 234567890Y� �f�@����?�W�( АP��8�h�х�ڎ���HR5ǃ��	��R�570�B�Aff ފ������ڟ�ǟ �"���F�X�3�|����i���į!�CE_R�IA_I�������F��;�Я ����GP 1.���s�H����V�C󠸾��Z��CO�C ��(��VǀC8��@��H��fCCX����Ch���p��x���� C�����Ⱥ��+�`=�G��ށ��HE/p�ONFIG=�f�G_PRI 1�B�$r�����������(�~�CHKP7AUS�� 1���� ,wuj�|ߎߠ� ������������0� B�T�f�x����DҍO���T��_�MORGRP 2�?� �\�� 	 �,��P�>�t�b���5�����e�.�I?a�a�����K����d�P�V��a�-`�/A�

s��������b&�i��ܦPD�B�����)
m�c:cpmidb�g��:�  C._+���p��U   � G >s��6� X��d�/�
/�a{C�e�/�./�/{g�+/���i{f/s/i��u/�
DEF ̋(K�)�b buf.txt�/�/���_MC������d,53����|ʇ�Cz  B��p�B�Z�B�X��B��~C� �Cޢ�D3��u
q�Dv��D�:�"Df��E�NNEA7E�V�ߓ=F�pg�F=C�Fi�W�G���Gp��OG�/�	ބ	6:����4���U(D~���/�	�ʄ3@à1
 TB��D�V@a  E�I�5� F*�� F�G$ˀF�[� GR�kNG�l��G��G���&H��G?֓�H��߃]���  >�33 ��ށ�  n4^��@߂5Y�Ed���A��=L��?<#�
 ���_�*2RSMOF�S��.^�9T1>��DE ��l� 
 Q�;�P � 0_*_>TES�T�"__��R�(��#o^6C@A�KY�B�Qo2I��B�0��� �C�qeT��pFPROG �%�S�o�gI�qR�u����dKEY_TOBL  6��y�� �	
��� !"#$%&'�()*+,-./�01��:;<=>�?@ABC� GH�IJKLMNOP�QRSTUVWX�YZ[\]^_`�abcdefgh�ijklmnop�qrstuvwx�yz{|}~�����������������������������������������������������������������������������q��͓���������������������������������耇����������������������Eъ`LCK��l���`�`STAT��c_AUTO_�DO��O�IN?DT_ENB;���1R�QY�K�T2�����STO�~��TR�L�`LETE��ފ_SCREEN� jkc�sc 	�UπMMENU 1i?  <�l�o l�K�u���FS���� 柽�ϟ���R�)� ;�a���q���Я���� �ݯ��N�%�7��� [�m�������ɿ�ٿ �8��!�n�E�W�}� �ύϟ�������"��� �1�j�A�Sߠ�w߉� �߭߿�������T� +�=��a�s����� �������>��'�M� ��]�o����������� ��:#p)+�_MANUALӏގ�DBCOu�RI�G�$�DBNUM�LIM�,1e
��PXWORK 1k�_-<_pN`r�TB_�  m��Y0�__AWAY��1�G�@b=�P�_A!L� =���YҀ��t`�_�  1!�[_ , 

:�&d2/o/�&�Mt�I�ZP�@P�#ONT�IM��d��&�
�e#MOT�NEND�o$RECORD 1'kqU2)?�!�O�?1 -?&k�k?}?�?�?88 �?�???�?c?O*O<O �?�?rO�?�OO�O�O �O�O�O_�O8_�O\_ n_�_�__�_%_�_I_ �_o"o4o�_Xo�_|o �_�o�o�o�oEo�oio �oBTfx�o� �/����� >�)�7�t�� pu��� ��-��͏ۏ����� N�`�Ϗ��o����)� ;������8���\� ˟ݟ����;�Q�گI� ��m��4�F�X���TOLERENC��B�	"�L���� CS_CFG �( +x'dM�C:\��L%04�d.CSVY� clֿx#A ��CH�z _/x.�G���},��RC_OUT )�- z/��?SGN *��"���#�17�-JUL-25 �20:52��27-MAY���14:38�]�? Z�t������x.����pa�m�?�PJP��k��VERSION ���V2.�0.11~+EFLOGIC 1+�/ 	d�������p�PROG_�ENB�2��UL�S�' �p�_WRSTJN� ��"��EMO_OPT?_SL ?	�]��
 	R57Y5x#?�74D�6E�7E�50i�d�o�2�E�d��j�"�TO � .����k�V_V� EX�d�% �PATH A�ʇA\��M�_�~+IkCT�F�, '��`�eg���}�STBF_TTS�(�	��Eм`�:��� MAU���.�"MSW��- )��Q},t���.�!�� ]l�R�v������4SBL_FAULy�/��#�GPMSK�ߧ"TDIA��0����`����!1234567890xS�l�P����� //%/7/I/[/m//��/�/�/�/�/L0PV ��� /�2?X?j?|?�?�? �?�?�?�?�?OO0O�BOTOfO8<x�UMP�$�I� �ATRp>�O�@PME��~�OY_TEMP��È�3��4��D�UNI	�w�YN_?BRK 1��x��EMGDI_ST�A	��_�LPNC2_SCR 27[��_�_�_�_�&�_��_o o2or�nSUQ13y_+?|o�o�o�otlRTd47[�Q� �o�o���_>Pbt �������� �(�:�L�^�p����� �� ?Ǐُ�0�,p� �+�=�O�a�s����� ����͟ߟ���'� 9�K�]�o��������� ɯ�����#�5�G� Y�k�}�������ſ׿ �����1�C�U�g� yϋϝ�ׯ�������� 	��-�?�Q�c�u߇� �߽߫��������� )�;�M�_�q��ϧ� ����������%�7� I�[�m���������� ������!3EW ��{������ �/ASew �������/ /+/=/wa/s/�/�/ �/�/�/�/�/??'? 9?K?]?o?�?�?�?�? �?�?�?�?OK/5OGO YOkO}O�O�O�O�O�O �O�O__1_C_U_g_�y_�_�_�_�gETM�ODE 15'E]fa t|��_GgRROR_P�ROG %�Z%����HogTABL/E  �[1O�o��o�o�ZRRSEV�_NUM �R  ��Q�`a�_AUTO_EN�B  u�SZd_;NO�a 6�[�Q}�b  *�6p��6p�6p�6p�`+�5pOastHIS��cXa�P{_ALMw 17�[ ���6|6`+t�� �&�8�J�x_�bp  �[4q�R����PTCP_VER� !�Z!6oZ�$�EXTLOG_R�EQ�v�y�S�IZ�܄TOL � XaDz�r��=#�
ނ_BW�Do�%��fQ���_D�I?� 8'E�t�TXa b[�STE�Pg�y��P��OP_�DO�v$v`FE�ATURE 9�'EQ��QH�andlingT�ool � DE�R Engl�ish Dict�ionary�7� (RAA �Vis"� Mas�ter���
T�E0�nalog �I/O��p1�
0�uto So�ftware U�pdateb� "�/�k�matic �Backup
�d�
!��gr�ound Edi�tB�  25L�CamerazT�FX� "Lo���ellT��L, �P��omm9�sh�ۡ�h600��c9ou���uct��p��pane� DI�F���tyle �selectѡ-� /�Con��9�o�nitor��H�d�tr�Reli�abT�ϣ(R-�Diagnos���Q�	�H�Dual� Check S�afety UI�Fc�Enhanc�ed Rob S�erv��q ��v	ԸUser sFr���T_i��xt. DIO Vf�fi�� )�\�wendܰErru�=L��  prנ*��rO�� @���EN�FCTN M�enuİv����.�fd`�TP In�?�faco�  
�E�G��p;�k E�xcذg�C��High-Speܰ�Ski��  Pa�r+�H���mmuwnic��ons��7\ap��urf�?�~X�t\h8U�^��connZ�2Т{ !�Incr���str)�8��M-�6�KAREL �Cmd. L��u�a��}��B�Runw-Ti�Env��(<�@�I�<�+��s���S/W�"H��License̾��� ad���ogBook(Sy>��m)	���"M�ACROs,��/_Offse\�f��b��H�!�Y�M1��MechStop� ProtZ�3� �5
�Mi4�S�hif\��B6S�MixܰQ�����H�Mode SwoitchY�Mok�*��.�� ��Mt�Q��g�� �5��ulti-T������)��Posj�Regi�>���  ! �P>A�t Fun1���6iB/��R�Nu!m�Y�3�G�P/��>� Adju��	��/2HS�)� o<(�8�tatu���wAD ��RDMޱ�ot�scove&� #e�v�㱗���uest 867�.��o�\���SNPX b��Y���)��Libr%�
�rt I���� "�����.S�o� ��s i?n VCCM����� j���������/I�� 710~�TMILIBXp����g�Acc��C/2�TPTyX�� �Teln���Y@����K�PC�Unexcep�tܰmotn�� �������\m725����w�5����  h640SP CSXC�i � xj*�� RIN��sWe���50,��vrl�زmenX" ��fiP-�a��x�P��Grid{��play F O`/��? ��ELR;��|�20��ORD�K�sciiw�lo�ad�41d�st��Patd��CyqcT�h���oriɰz:�7c Data� qu6�2�0�*��������FRLa�mc�K�HMI D�e��(����k�PC��φ�Passwo�rd�644��S�p�����D#YEL?LOW BO�	?1��Arc%�vishu����#ti�Op��^�! 2��aO�p�o�� t��ֶT1�o�����HT��xyy�	�   $�t۠ig��10Ơ� 41\+�JPN� ARCPSU �PR+�8b!OL�0Sup�2fil�� �!��E@-�;�croc�82��v���$� 12jSS0e.4�tex-� I�7��So��tf�ssaEg�� e��У�P���,��� "Tc Vi#rt��v�!����gdpn�
�J3��SHADf0MOV�E T�MOS �O TԠge�t_var fails l�>PU~1�E���� Hold_ Bus %�h���VIS UPDA�TE IRTORCHMA A�{�vY�WELDTV S �]�DtS: R74-1��ouiPb}�y���BACKGRO�UND EDIT� "RC$REPTC�D CAN CR�ASH FRVR� 62z1�SCra���s 2-D��r� ) "��$FN�O NOT RE���RED �` m� ��JO� QU�ICKaPOP FLEN m41S��Loc��gRTIM�Q%�#�FPLN:� FG��pl m�r�`�MD DEVI�CE ASSER�T WIT PC�V;PB�AN#aAC�CESS M .�pc��Jo��Quqi±�Kbldmg�USB$ ��t &� remov�� �Pg�SMB NUqL� ;a|�FIX��}C��ACHIN,Q�OL�`MO OP�T ՠa��PPO�ST0�WDU C��wQAdd�`ad����0io�2��$�P�`W\0.$0`O��IN&�P:fi�x CPMO-0�46 issue�C�J/aO-�0�r1�30Т- ��vRS�ET VARIA�BLES-P{��R3�D m��view� d��M��&�ea����b��of F�D�5P:N@x O�S-1y0`�h s�c���t��s t�l�o��7 WA�PZ�3 CNT0 T��/"�ImR�)�ca� �Pu��POT:oWhenapewB�OSTY E�{1t���ptKQdo GE�T_�p �p��VM�GR LOl�REAd0C~QW�~1�(�pl�s�gD�ECTp�LpING IM�PR�DR(p+PB�P�ROGRAM�ER�IPE:STAR{TU� AIN-;��ӠM/ASCII<zPÂOF Lq�DPTTB: N�p;ML$me P����`:x�mo&�alqlW`!�ӤTorc�!A�U�HC�iLpԸ�th�`n�@ ch��/GEA�!�tou<͐�RCal��k�oSign`� ND��ԗThresh1�23��`��09p :? MSG_P�+0Ger  �Q�Aܠ�zeron��0 gH85��RImA��n�2D��rc�0I���OMEa`�pON�aP5�  נSRE#G:FF-Д� ]�'����KANJI��nʖ�J��c�0asn yd�!OA immc ��INISITA?LIZATI�����~1wem����dr>+� LB A�UWq�minim�reAc[�c!�R���m$�ro -1>ѮS�ܰir��@ұJ�1pd�ETw�� 5`?�I�o�w u��< se W1lc��YbPM����p�Q���R`vR&�lyu\�3�Re 0�d4q�q1#���m <a��arn��ঁB�ox fo��*PR'WRI�PW�S��v�k09 F�pupᐿde-rel2 d��p� j��`━be�twe��IND �Q���igE sn�ap|�us��sp�o TME��TP�D#�DO�p#aHANDL 1\k�`(vR��ȀD�ny�S��v�Yoperab�il� �T*�: H$ � l\p��Vq�b��R�< p�a*�c&2OƝ`FA,�.�-QV7�. f.v��GT�pi�s��� ɠ�tmLine-?Remark ��/ RM-�` W�#SPATH SA+P�LOOS UIF�c�+5f fig�pG#LA����Vrp����z��U�0ther�>V� Trac���tW�\b�s7��d�ht�� n�@  ��R�3:���dK�y���it k8�d�Pa�yR![2]�ü1�: g��s��doew�XQ��0IS�q��qEMCHK E�XCE C���M�F +�Xah�� 35\k��)���QBt���'b���[�c���e �`k�S�� BUGr��cD$`PETp����f�c4��0XPAN;SI��DIG��@�OoPmetTCCR�G EN��CEM�ENT�A M̀K� {�`H GUN�CHG �`� EX�T�P�2�bQS�9�3 wP8�x�ORY�LEAKq  H�5gyq�PLC W�RDN R �O �/u�QSPE=p��G*�V ��$�tn7w20\3pGRI���A�rT�PMC gETH��pSU7p��`  j5/n�PENS�PN,��*P� ont�`BRO�W�`!sRMV A�DDz CN qD�C���PT3 AL�A2@ ���pSVGN EARLY�R��ŰH57�Ga�JLAYҀE (�@M�PPD�p*@HΐS I`P�OU#CH8���V�F�q��comH�x ��ER�ROR� DE n�J��RO�CUR)S8pI��N4q��-158n7�R'SR xP#aUp��(�Rqy�T�Fz�;`�pk��t�� gՂ��B�SY RU;NN�  a�`��BRKCT�!RO<�p3@ \apSТ�cAXxP���h8+ <q��ISSUr} �sPX�PTSI�K�1M10_�IPSAFETY Ck�ECK[��Á�������<#X�� �TW�D2�@�@�INV���D ZOp�5Xx��t�DUALy�� "M6�0�"rF�#�E��dPdNDEX F�t*UF�"Pʀ�0sF�RVO117 A��PT6�KtqFAL�PTP2477D6r_�P�!;HIG� �CC�t;SNPX� MM��tq�d~ҁVq�q#�
"��DETEC�Tq*@RRU�qA�P�5p�9� y�)<9���7T���Pds� k��	���!Q���� �t\4A�;A0�2 "Ke@" 8@HI�q�XF8@4@H�PRDC"�
�aMB8@�IXF�b���zOX@8@���a�G}E�B�Ccscr��J8@�Ndctrl�d.�A�NZE�A5�$�Q��!�`�Df8@�`�m�878�Q-;� ^��� rm`�
���PR̠78�@RI08@0q�Q (~\Mp@��0t��!{B8@\tQ�<OX�St0�3hB3�nO�Vtp�A�@LC�F�L��� �Rpl�cf���J8@�WTam�ai�E8@mubov 2_miTA�O�S8@U`T[xtT�AqPr674xS�Shape GeQn��8@j�I�[R�`ĝ@8@T����%q (u8@��II�^�Q~C`�a�[8@;Ynrsg0��4� � 4�CtMr)68@�r5hB5�zVnnretsp "r��Po�wng0bGC�RE�Ka�ޠ�D�AT�E�k�creGat.�q�M�a�o|ksqgtpad1P<��(�tputZj�{ �������܆28@��0��Q����sl�o��;� �hexH�TBp�8�ď�keyH��8@�pmZb�NR�u7A+�nrgc8@UQ��pp�bUZ�dp0aj9�21xSpl.Co�llأcq�\A��RN�q�UA� (J�8@ip�_�WA��_�Y��ae7hB7�ͦtp[�? "TCLS9oKb��clskyh[��s�pkckZd����$�TQ���dA�rx�7�10a- KARE�L Use Sp��FCTN9�a�70l�0s0a�� (���a���~C8@��MI��c8�hB8"   ��8@ v	��v	   lm7atea99�qM�����E�mcclm5�CLM;�� �j��fE�et���aLM	��h�yasp,���mc_mot�B�N��8@0H����Q��su'��Q��ȕ�䅮���joi�#�ߕ��A_log8�Z���trc�B����ve�ϓ�v��QWX���6�finder�xSCenter qF1�lSw520���ha6rX� (<�r,�Q�Ձfi�Q �NH 0�I�ۡ���A8@uL���tq�a "FND�RVϳ���etgu;id�UID�C8@����������TA@�nuf;��P���ƞC�B��_z�Ӡo��qG�������l���fnd�rTY��2䁴tcp<"�,qCP MF�}�38@517��6s38�E��gf6��(� �K��Q��-�X��A�tm6�P�İ� �Q���	�͘��Ctm�Ĵ�b8@ej��TAiex��aP�Apa�ذ�cprm�A���l�_vars ��
��dwc7 TS���/�6��ma7AF�G�roup| sk ExchangJ �8@�VMASK H�5�0H593 H�0aH5@� 6� 5�8�!9�!8\�!4�!2���"(�/��;OMI� `@a0hB0`�ՁU4U1#SK(�x2�Q�0I�h��)�m�q�bWzR�Dis�playImQ@v�J40�Q8aJ�!(�P��;� 0a��0���� 40;�qvl? "DQVL�D���qvBXa`�uGHq�O|sC��avrdq�O�xEsim�K40sJ#st]��uDdX@TRgOyB�Bv40)�wA~����E�Easy N�ormal Ut�il(in�K�1?1 J553m�0bD2v�Q(lV40xU)��������k986�#8Uϕ�|�rP "NOR��dw d.a}oKksu�O�W���OY��W`�j0�6�H� me'nuuyP6�M�`wR�X�R577V�90� �RJ989}�4�9b\�`(�fity�����e�<?��&Vsmh`��8��C0�Sv�q�8���w��pn "MHMN <��ޣx�Ay`�o�3�u �`f�І�x�t��t�RzQ��LV��vP�tm����|I�1{oPx �2�|���I�3I/B�od3stǏًmn���^�}ensu_�L<����h!!��Rt��huserp��0Ҹ�ʐcM�_l�xP�oe�<�рpoper���>�xdetbo/�l> �x���Ps$p�`����OPydspweb ͓��z'R��u�Rr�101&S՟{t�`2�Z4�30�����"�`4�
�4�5��KQp�m[T��dUCalG 40`�Q)p40}������9;��DA�� �v	LATAum�pd�\bbk96M8��68c�fbl�.41969y�9�|�D����bd� "BB�OXêM��sch�ed����m�setauM:�����ff� ��40��n�41�ϒ�40�q�col��|�1�x1c�ؘ���li��X� 0���j��&�8�4 <�{ro5�TP E�l#��ryK42r���;�(T+Q �Rec'�ʈ1Iw�84��x���Ak971���71�;���parecjo��QNS��[T���dXrail| nagek�M ,QjT2 *� (�ĜR%<x�80!bTh��p��4��4�y�Dgl�paxrmr "XRM�g�l��brf{���n��k�l��9turbsp���㧑- �l015	�g�625C�Mh� +���)89��	+��B6��o�ҹ��x��7�q40����pd? "TSPD�=��tsgl��l�:`dQ���8Bct���K�vrE�aܮ������  1�!���21�`( AAVM �2��0 �@fd T�UP him (�J545 ly)�`8 616 %�VCAM ��CLIO (��0:�5&  (=F\ MSC �Rt"�PBsSTYL��D!28 :2\ N�RE F2h SCH�6pDCSU� tpsh �ORSR �rD!0�4�SEIOC�& \fxh 542� LEX"� ES�ETn�8!H ��sh�8 7H �MA�SK�Ø"7>��OKCO*`x�!03"6(�!/400:66$ G6s39.6[8LCH!6oOPLGR703
5OMHCR��0C� h(! �06�A.f8!�54
��00DSWb 588�180 �h!�37 88 (D��"02C24���27 q9�25��2-6��05��9PR�ST bBFR�DMES�!zB�9�30 _ NBA�  6� HLB �3 (~!SM�@ �Con� SPVC� �8!20z��T�CP aram\TMIL A���@PACETPT�X �@p TELON 96��29�%�UECK��r U?FRM et�P!�OR ORP IPL^%CSXC�0j�1�CVVF l F�QHTTP st�A")�I#� CGHP8~ZIGUI�0��hPPGS To�ol� H8�@dj`Z��!@�h!63�%j�@32Q\�31 B��h!96�%R651��Rs�!53 TF�AD�R41�8"1� ��oo�"9��41775�"/@�P�VCTO�@�U�!sh!{80�%PRXY�R��!770 �b8 8�85 ol3P� L� аdi� �`ڳh �LCP{Q� TSS� �b�26:����@C�PE �HT@VRqC~�tQNL ��@002 %��b	0gdis� �`7 <°�a\0�T�`1 �`e=n�b4 652�`)FU02Q0Πo`p2�Ptu�r4 $r�5N��RU0p@ns�e�QJp1 APFiI[ Jp3�g34�g40 alxrE1�t44w46� ts U0  7v�0O��r5�e�p7 p 7"sw�a61:��rY4��r5 QpwGr�`�$�p8R�"sP`tjQ�b�36w77�wL8`�v83���r8�&�:��pOq8�8 "r�key8�9F��a90�91 p�#@���� �D095�g97*pur�A1@d��H�P|P�q1�0QplSqA1p#4��]a!s1@sl༂8�Ӽ�\1�d1�`��v�@{��14p�ae��5 hH2��`�6ޣ��7�f1p@��d�YpCqd�ـ
d�1�`uq��� Cu�1< Oq� ��7ReU	1$ �u1�Pϱ� ���@- WQ158� ase C��9� B��60 82�ń�p���4 (W�ai��`吢!��7�E��8�EU1P`rIo9�<�1��<�2��<�	0��T��l�5HJ�l��cC���9%�GMCR��P�2�`t�Q2@967�QR��8��9Z�2TP�B���P�2P7U5 @�o���
�5�`U���3 w���?A�E$�1��c�qAwl��A��1��512 f���1�u5Р���a5p$��56�+a��Q15h��Ұ�1 @���pp�b[�538 BxaB��|p�4�2�1e1/q5�p�4U5�P16 (߲�Pz��0��8�P�����p�e5`�e5(�/�P`bbf>�X��$Z�U�}5d�\� X¿7 	  ��8� k_kv��79� s�82 &�H�5��E6���p����h ���ñ���3J"�`n��4 3Ȥ59ѧ�6�0t���8��6�D0$�$�4 7���!���<�j670\tchk<�Ps��<�B<�90��7�<�$��<�\K�<�q�Ӻ� A�C<���q�<���<�mt��sg<�lc���FA<�H��<���0<Я���<�hk��<� ��B<е�o�<���<�x�K�<�dflr��<Ш��� ��o�`����D�;�<�gEvam����B<г�oќ����<а�KЀ�creexl����P��<�X��|���j6<�s��prs.`���\����<�7������fs�gn��P�b�t�at ��<�L��1B !��svsch/  �S�ervo S��usle>�SVS��44�1u�_<��� y(����ched���,��~��A\��  �� B���B�qA����Zcj�� � 5��1<���Ә�p�cs?s "ACS<�& (��6� �����c el���Q����?torchms�<�7- T�Ma`Ѵ���09 J5;598 J681s�7� 8��b��<�p�a����te,s������/�E�� �m��ARC.�� 1q�4�!=��C�tc�pA�@t��Ѧf� F����7#�2x�SE�r���UstmS�0960'���RC����0��� p��96G= '��"H5W����L���\f�� �@PATb���`!4U�#!Stmt�E `��� �pMA�!�p��z�2?�in_�<�X��r�X e/c�W����V����e�tdl�vߏ\ov�eto���܏��m?monitr�\��|#�0st��?.6�a��PP���!� Q�!y`�`ame� �Arol�c�43�0 �p��ћ01� 25� � �<� v�	�v	�A@�818\n; <s�I��B�2�pMPTP"���C�1mocol ��,��CT�v�'!� �A����8P53��y`T/ouchs�s�`��<��J5���Ѩ`mP����n[PQ�a ,�E�a��IP&
�Pth�A<�KF#R�m;ޱQetth�TH�SR'�q-�Rt��o? "PGIO�#!$�s�ISwka�"WK���!�MHqH5�4��5w5n/�Sm/��@ 7�*�da���8`!w/Ac��tsnf Tk�/�#gb�aP��u`��^m�`u��Zӭ�ܱQp�є�#����Ka<��M��t5 QtZ�a<��dFS5GhK����G�1or��dW��64��tPx���P ����x,��?�$���P<�Z4e7�g? "SVGN.ox��copy "CO�;�Wj$�O�A�9� "FSG�ѧ�%7��_j��f� wQSWF*|!"(�sgatuɀ����_
��tp_T�PDo��9�79��#dߎ?���h�GA�T���!#��  �Гf�` ��"/� �w�Z� �b?6?� � ���� ���E ���M� �chrT� �K6K� �sms� �o6�ѐ�?gtdmen?3 ��?��� ���mkpd�td2 ���, ���pdQ�X� ����� ���mvbkup. ��[�C�С��mkun�o��prp���mk�l �4��s �nixU��� �ldvrw���glg�4�� ��渣���aut7�.pб�旐 �ַ������su3� �Ǜ� ��Ƿ� ���\ �6�b2X� ��&�� ������A4�  ��B   946" ���fB� �t\pai�c\p4k947� ���F#���� �icgtas���pa`���cc:�<��o���N��gen�� � �F�lnp � ����sctf@��1��wbO��c��Ջ�`��߄�vri�ߢ�а�-T� �x��p�flow� 6OPAc��ow���R50qtS �#T� (A��4�#���p��V�cu3�QF� �̾SI�ac����46`����s&��pa��`!!���� ���55�b  �o)�p���0娿
��afcal3�P� @��f��}���`�f��m	߳�p�d�m�/���a/��$C`ѷ�� �! track\P�� 0�ine/Rail Tr�]TJ�s69W�T  (L�� 8(`љT.�`�%��HD��P0� (��8��48��_ɛ�⇒4������ �3�b3����alV@ �N�Tf���%��Iinp]0m���aen�� ����&?5�c@Itst3@��$�� ��`�,R9�%���0�氱%��pope/ners-OW dGDev��F�M�6W����|A�Pc"�l!esv� �,��R��V$�Q`���U<�V$ �k9j 
�6��# �����%�paop/!OPN�U�V ��2celL��8g_��/�6��tscG��$��V!��3� 5vrop�ߡ�7`�n(`�V" 2D�a V'O$:S9�>�� PumpE�� jQ�@�" ��!
��@бMSC#�@��)P��AC��`��� � v����� \mhplug�@g�"7P���uK")㠱io7�CpJ0��E�LIO q51g 7A93շ�E5 q9 t����4rb� ST��R��CPJ�989�P�LSE(�' �e C3Q(P �/Ov���o�P�� ? I1�R���55���f�I1`�tcmio��MIO�����U�tco1"CL01dV �cBK`io��uM?���Sl�I0�߈��Eg �o���f �tI4\onfdtI����e%�p27�Inte\�TB CoMoo1�E�R�(do55G4 (;r>Ex,�8�nR##ipc�/>�&�qp5���
oQé�1�p����7/o���r5a�pd�CDV_���rP�֮��qp2cnQd��s �p��a�o��r`҄�S��"�c�a�c���2kIԿ?A�pcrt���or0�qd#��"���3p+����D��Џ��vr2k �0���AG�.+��gcho�;�uC��8(� �uV630�fw e P�mී�@���`���TX�� ��d�chp "_��(	��3�����8����\p3�v����ш�9��3�1 �����laow�[ͧ���chk���㳦s��s?Ө0�i�1h���2��i�w����s?1*�-	�:�O��vr������p0�'���PFRAPwWat?1rneE� P�sp�& ac5� _A.�rbo#�,�a��g��������Qs<�ICSP+ 9�_����� ���F�A9PH51IQ9%3 7��HX6hQ]PdVR`S5��fPR6 liQWPR� (P!/am S�u�"�A|�I0�tpprg�0���`h�@2atk932�!��E�^��a/sc "8�C��S>i�atp�"�d�@1�I�
g�dsbl�fltJA�Qsab?le Fau�P{�C!��EV0ex/!D�SB (DC��t �$�p��X 7� �� 5��Q�t3*�~��6��td9� "!%�(5��sb9኏����\	�6#���@5�p$�D@550-Adj�ust Poin	tO"tVJ�Rs�z�� ���!�X_�Yj��/0\sg��4��}7�y�\ada�"A�DJ���j�Qet�sha<�SHAP8�sŭ'jpo�r4� t�!��$ ��C|��	Tk!bRPKA�R/Qiagnos�tì!O!vV66C J`ew0�(��L���/�&krlde� ��PP���hUH b���r3�Pp?q���DBG2C��� ��X�o�1U�� `��WT`�@ipJC�M�aipper �Opv`1Se}78? (MH GF�  ;":�&##�� a�x��,�$��388C���(��#��9.�9C��g$##PPk�Q��8�!�_ "$�"��=0%�P��A $���_�#%0AQ�C~2 �Mat.Hand�lE��!= &�pq M�PLGET�0�1( �3�Tt&P�Sٰ'�B� 1��B0����&p��H�� PP �'p��@�C7PP@	�TG�tD5�}m�q��Afhnd "F~_R  �����>PP	   xT?Qܣ��P(Pa��To������?�pmpa�O��JP ak925B��2`@O�JRpsQ�`B2�unLHP�Tgse�GSo1�O�W��QT��v !�R�Pt�p~���JRdmon0.�@��V�!ns�hYvr�QJ�g�Q�o�jXY�HS~7sl�f ��pen�PDnR(R&���ɐ823'��ٔ q���g� ���� 1��� S�� ? �c\sl tQ�!|QE�P��a�rtP�g��P�� �v��"S�EDG8�s0�qtdgY T����v P`ho�s`<`����qc�`g
�e` o�w8�a@o"�ile6�H�e�ȅnR�� �e<! j517�>����J%��e�`��BQ4��Q&�L�!F�J�=�o�5�z/l17���_�œ��`C�0C�  ���LANG j��A��������gad���,#�jp�.��4�Ē�ib���s�Ƒpa���&�~��j539.f��,Ru� Env�
������3H�z�J9�����h�Ф
Ҕ���2�2����� (KL�n-TimФ�⠤���p�3�TS����\k}l�UTIL"o����x�r "QMG�l��!������1 �"��S�T3�\kcmno��SФT2�椱ut�.�lre3adc�}�exY�ܤ�r��\��l��Фw�a3��2C�*� -� C�D�E!Ĥ� .��C�� R CV̴�Ҁ�\�p�Р���p�t�box��.�@�cyscsL�:�RBTE��veriOP�TNE���;ӕ�k�e`�ߦ�a�ߦ�hg����DPN��gp.�v��r�ptli�t��0�4��te�\cy����tmnu3`�r���5UPDT��������駣��it�e �� swtox�,���oolB� F"�Y���Q��(q��gr3��䪒��"�䂴�w������߳��s �������������ylS���bx "O�� ����l����P���A�l\t�� ��p������	�Col�9e!��R C��r���&r �m;`��Chang�Lq�T1 �rcm3�"��
� A6���"����sP7���"��222���2D45�7�� CCFM��H��accda��Q�c' ��KÕ 0���K!����mo!�� �,$Á��!"
� ���/�/����	Y�,$0��)�,$sk����
m rC%tS1,$+��<k1�%unc.,$o�8��1��sub����8��1��cce�5/�!&��-/?-W/i&v s�}/�%#�#�/�.C� �/� C%
�@? U �&�+��F:qt�
pD��� D	  �U�:7�Dxmov.�P��DPvc5Q�tfr@PeC_UYg�eobdtg_y[tAu���P���PTUt�P��Sx�_�^z�_�\v3ar�_�\xy�_�[pcl`c�P���P��Ue�Pgrips9uaoskuti���o>vfinfpo}��o��j�b�P���Qud\@�aX��Pc�\Rrp�QAnƅ�P�v�P)tm#q`Ɔ�P�v�a+rog�aࣆ\Q�?a+rpal?a{�{spa���P�u�Q�t�_TZp�0�osi�pkag3r�ovlclay(�:�t�p�T�d�pu?a�c�A� �����KtKa�P����9qTf|rdm��{Grin#r���s� �2���|s�Pd�v�tv��v�h�0��yGstn* џ�yt'�	1�p��D�p�uϑ#�Cul�@o�W6�2��siupdl�]�o�vr�on��`1L�z�`8\�r���il3$|#l4��ǉ#q54Fy�B�Տg{�`���{wc�mס���wxfer��UYtlk2pp<߿UYconv��si�cnv�Qʯxag8��H�Z�lct`ao��=�p��׭nit0�믁�3������  ��� v	��v	$��alFϑpm�r&�B�eWa ���f�%�������I��߬�u�ͬ�Kam�T�f���c��w��ro�ǁ#�5�����?� sm ��y�a��y넑�� ����`����͐ϑ��p��m�Wa�1�� �A�6�S�e�X��ψ� \Q}�����������ĥ w߉�西߭���߮� #q0��rs�ew��� 1�a��z긱n@�.��۲;�d�������  � Ad�	T$�1 p!� P��e �e �	lf@C�@��s/�  ?�����8� ��������reg�.�C=��o9�9 ~@�����$FEAT_IN�DEX  z ���e�� ILECOMP :���1!�!z$#S�ETUP2 ;�1%;"�  �N f!$#_AP2�BCK 1<1)  �)��/�/G  %�/�/e4  �/�/>%�/$?�/H?�/ U?~??�?1?�?�?g? �?�? O2O�?VO�?zO �OO�O?O�OcO�O
_ �O._�OR_d_�O�__ �_�_M_�_q_oo�_ <o�_`o�_mo�o%o�o Io�o�oo�o8J �on�o��3�W �{�"��F��j� |����/�ď֏e��� ���0���T��x�� ����=�ҟa������ ,���P�b�񟆯��� ��K��o�����:� ɯ^�����#���G� ܿ�}�ϡ�6�H�׿ l�����ϝ���@)t �Px/ 2� *�.VR��߅�*��@߂�F�j�T��P�Crߛ߅�FR6�:����V���z�T  �!���K� ��<q�S�*.Fߢ�"��	�Ӑ���^�����STM ��'����S���iP�endant POanelS���HI����9���U�������GIF0;��������JPG��;��]oR�
AR�GNAME.DTy�>�\"����Rc	PANgEL1Y�%>� ��e�w��2�A/@�//���/�3_/��/��/p/�/?�4 �/I?�7?�/?�?�TPEINS.X3ML�?>:\�?t?��1Custom Toolbar�?�Q�PASSWO�RDg?w�FRS�:\:O�? %P�assword ?Config{OR� �OSO�O�O��_�OB_ T_�Ox__�_�_=_�_ a_�_�_�_,o�_Po�_ Io�oo�o9o�o�ooo �o(:�o^�o� #�G�k�� �6��Z�l����� ��ƏU��y������ D�ӏh���a���-� Q���������@�R� �v����)�;�Я_� �����*���N�ݯr� �����7�̿޿m�� ��&ϵ�ǿ\�뿀�� y϶�E���i���ߟ� 4���X�j��ώ�߲� A�S���w����B� ��f��ߊ��+���O� ��������>����� t����'�����]��� ��(��L��p� �5�Yk � $�Z�~� �C�g�/�2/ �V/���//�/?/ �/�/u/
?�/.?@?�/ d?�/�?�?)?�?M?�? q?�?O�?<O�?5OrO O�O%O�O�O[O�OO _&_�OJ_�On_�O_ �_3_�_W_�_�_�_"o �_FoXo�_|oo�o�o��`�$FILE_�DGBCK 1<����`��� ( �)�
SUMMARY�.DG�oblMD�:�o*n`Di�ag Summa�ry+8j
CONSLOG qn��=qConso?le log�7k�pMEMCHECCK��2��q�Memory D�ata3�;g� {�)�HADOW�(�����C�Sh�adow Cha�nges���c-��)	FTP������=��qmment TBD;��;g0<�)ET?HERNET0�`n��q~���=qEth�ernet �pf�iguratio�n��B`%�DCSV�RF/��'�@�C��%� veri?fy allC��c�1p� �DIF�F8��0�ůD�%=Z�diffǯ{���q�1������J�c X�q�|�	�CHGD�&�8�ͿBD�ܯ�����2Ŀ8����R� `�y���GD�.�@���D�q����FY3��8����Z� hρ���GD$�6�H���D������UPDATES.$�
�ck?FRS:\"�c��>qUpdate?s Listc�`{�PSRBWLD.CM��blN��e���pPS_ROBOWEL\�6o+�=�lo a��o����&���J��� n�����9��Jo ���"��X�| #�G�k�d �0�T���/ �C/U/�y//�/�/ >/�/b/�/�/�/-?�/ Q?�/b?�??�?:?�? �?p?O�?)O;O�?_O �?�OO|O�OHO�OlO �O_�O7_�O[_m_�O �_ _�_�_V_�_z_o �_oEo�_io�_zo�o .o�oRo�o�o�o�o AS�ow�*� �`���+��O� �s������8�͏ߏ n����'��� �]�� �������F�۟j��� ���5�ğY�k����� ���B����x������C�үg�v��$FoILE_N�PR]����Y�������MDO?NLY 1<��U�? 
 ��ۿ (���L��5���Y�� }Ϗ�ϳ�B�����x� ߜ�1�C���g��ϋ� ߘ���P���t�	�� ��?���c�u���(� ����^�������$� M���q� �����6��� Z�����%��I[ ���2����?VISBCK����>ų*.VD�*>� FR:\V�� Visio�n VD fileVd����� ��	/./�R/�v/ �//�/;/�/_/q/? �/*?<?�/`?�/�?? �?�?I?�?m?OO�? 8O�?\O�?�?�O!O�O �O�O�O{O_�O!_F_ �Oj_�O�_�_/_�_S_��_w_�_o~�MR_�GRP 1=���LeC4  B�`	 ��lo~l�i`۬B���D��fn���MT� ��� ����e`i`a �o�khb�h�o�dc�ic.O�V�L�PK��t�M�SHIʇE��|�i`?���"B��A�f? �BO�9���l}�A�fA���A�ψAݼv�A���pl}F�@ �qhq�y�~g��fF6�D��MqD�� BT?��@��Ô~p�D��6���l����5��5���|�l}BiHZ�B��`B�$��B4�Bg���BWqr�~e9��BhFaA����A�}�BE>B�dl叐�A�����A�܏e��P���t�  @�C�m@PK_<`�>@�	Ƙ���� Ο��+��O�:�_����p�����eBH�` �����A�Mb���'�d
���Z��WZ� a�/�FX
�A@�~��@�33@���'�\��[���ѿ��@��񿋯�*���N�9�r�]ϖρ�<��G�=�<��m]<�+=~��m<c^��8�eN7��7�ѷ7�x7;��51���	ߤϨ�?߾d2^`Yb`�*b`�����F�`�U�b` b`�0�����C�^o�߂o�o �߸o��o�� ]�(� ��l���������� ��#��G�2�k�V�{� �������������� 1 ��-�) �������0 T?xc��� ����/')�'/ M/_/q/8��/�//�/ �/�/�/?#?
?G?2? k?V?�?z?�?�?�?�? �?O�?1OOUO@ORO �OvO�O�O�O�O��_ ��J����`_*�_N� �_�O�_�_�_�_oo 'oMo8oqo\o�o�o�o �o�o�o�o�o7" [Fjh�x� t��!��E�0�B� {�f�����Ï���ҏ ����A�,�e�,/�� �������/�J��� �=�$�a�H�Z����� ����߯ʯ���9� $�]�H���l�����ɿ ��ƿ���#��O�OV�  _z�D_V_��z_�Ϟ_ ���
�C�.�g�R� ��vߛ��߬�����	� ��-��Q�<�N��r� ���������)� �M�8�q�\������� ����������7" [Fk�|�|�� ��֟3�WB g�t����� /�///S/>/w/b/ �/�/�/�/�/�/�/? ?=?(?:?s?:�LϦ? p��?�Ϧ� O��$O�� T?]OHOZO�O~O�O�O �O�O�O�O_5_ _Y_ D_}_h_�_�_�_�_�_ �_�_o��@o
�go*o wo�o�o�o�o�o�o	 �o-*cN�r �������)� ;�M��������� ˏݏď��%��I� 4�F��j�����ǟ�� �֟��!��E�0�i� T���x���ï�?�?�� O��?OO�t�>O ������ѿ��ο�� +��O�:�s�^σϩ� ���ϸ������ �9� $�6�o�6o��Zo��R� ���������5� �Y� D�}�h�������� �����
�C�U��y� ����d�����:����� +Q8u`� ������ ;&_Jo��� ���//گ4/�� x�j/4��/X�n/|��/ ��/�/!??E?0?B? {?f?�?�?�?�?�?�? �?OOAO,OeOPO�O tO�O�O���O�O_�O +__O_:___�_p_�_ �_�_�_�_�_o oo Ko6oooZo�oZ��o�o �o�o��xo
G2 kR������ ���1��.�g�R� ��v�����ӏ���	� �-��Q�/*/��N/ ��r/�/ޟ�/��/)� D�M�8�q�\������� �����گ���7�"� [�F�k���|�����ٿ Ŀ���O�O�O��W�B� {�fϟϊ��Ϯ����� ����A�,�e�P߉� t߆߿ߪ��ߪo�� +�=�a��߅�p�� ���������� �9� $�]�H���l������� ��������#G2�W}h�p��$F�NO ������W
F0� �  #��1 D|�� R�M_CHKTYP�  � �q�� k�� ��OM� �_MIN� m���}�  X� �SSB_CFG �>� ~�Jl�Aj|��TP_DEF__OW  m��>�IRCOM� ���$GENOVRoD_DO���n�THR d��d�_ENB� ��RAVC_G�RP 1?3� X�e/��/�/�/ �/�/�/�/�/? ?=? $?6?s?Z?�?~?�?�? �?�?�?O'OOKO2O oO�OhO�O�O�O�O�O\�O�ROU? E�. q����>��8�?#�O_�_K_m_o_ꐖ  D3���_E�_q�@A��\Bȡ��R���>Y_6 SMT<#F�C-�Ufoxo�o�HoOSTC,1GYn?��_ 	�hM�k�o�f�oyeCUgy �z1�������p	anonymous�5�G�Y�k� w��o�o�o���� ��*�<��`�r��� ����ˏ	����� &�8������������� �ȯگ���M��4� F�X�j�����ݟ��Ŀ ֿ���I�[�m�ρ� fϵ��ϜϮ�����}� ����,�O�Pߟ�t� �ߘߪ߼���/�A� C�(�w�L�^�p��� �ϸ����������a� 6�H�Z�l�~������� ����9� 2D V��z������ #��
.@���� ����������� //g</N/`/r/�/ ����/�/�/?Q cu��/[?��?�? �?�?�?)/�?O"O4O FOi?�/�/�O�O�O�O�9m�aENT 1H�[ P!^O_  `_?_._c_ &_�_J_�_n_�_�_�_ o�_)o�_Mooqo4o �oXojo�o�o�o�o �o7�om0�T �x�����3� �W��{�>���b��� Տ���������A�� e�(�:���^���������QUICC0 �̟ޟ?��1@��.����2��l�~�߯�!ROUTER�௼�ί/�!PC�JOG0��!�192.168.�0.10	��GNA�ME !�J!�ROBOT���NS_CFG 1G�I� �A�uto-star�ted/4FTP:?�Q?SOBχ?f� xϊϜϮ��?������ �+�߿�P�b�t߆� ��6�����(�J�  �1�C�U�g�6ߋ�� ��������x�	��-� ?�Q�c� ?2?D?���� �����)��M _q����:�� �%t�����m ��������� �!/3/E/W/z{// �/�/�/�/�/6HZ  ?n/S?�w?�?�?�? �?�/�?�?OO<?=O �?aOsO�O�O�O�/
? ?.?0O_d?9_K_]_ o_�_PO�_�_�_�_�O �_�_#o5oGoYoko�O �O�O�O�_�o&_�o 1Cogy�� ��oT��	��-� |o�o�o�o����o�� Ϗ����)�;�M� _�q��������˟ݟ��ÿT_ERR �I�����PDU�SIZ  �^ڴ��$�>=�WR�D ?޵w�� � guest+�}�������ů�ׯ��SCD_GR�OUP 2J�� �`�1��!怒L_���  ���!�	 i-	��E���Q�E� EATSWIL�IBk�+��ST 4�@���1��L�FRS:�аTTP_AUT�H 1K�<!iPendan�������!K?AREL:*���	�KC�.�@���VISION �SET���u���! �ϣ��������	�߀P�'�9߆�]�o޽�C�TRL L���؃�
��F�FF9E3��u����DEFAULT���FANUC� Web Server��
��e�w� ��j�|��������WR_CONFI�G MY��X����IDL_�CPU_PC�惑B�x�6��BH��MIN'��;�GNR_IO�K����"��NPT_SI�M_DOl�v�T�PMODNTOL�l� ��_PRTY���6��OLNK 1N�ذ�� �2DVh��MASKTEk�s�w�Oñ�O_CFG��	U�O����CYCL�E���_ASG� 1O��ձ
  j+=Oas�� �����//r.�NUMJ� �J�� IPCH�x��RTRY_CN��n� ��SCRN_�UPDJ����$� �� �P�A��/����$J23_�DSP_EN~���p�� OBPROqC�#���	JOG��1Q� @��d?8�?� +S?� /?)3POSRE�?y�KANJI_B� Kl��3��#R������5�?�5CL_�LF�;"^/�0EYL_OGGIN� q���K1$��$LA�NGUAGE ,X�6�� vA��LG�"S�߀���J��x��i��@<𭬄�'0u8������MC:\RS?CH\00\��S@�N_DISP �T�t�w�K�I��L�OC��-�DzU�=�#�J�8@BOOK U	L0��d���d�d��PXY�_�_ �_�_�_ nmh%i��	kU�Yr�Uho�zoLRG_BUFF� 1V��|o2 s��o�R���oq��o�o #,YPb�� ���������(�U��D/0DCS �Xu] =��� "lao����ˏݏ�3�n�IO 1Y	# �/,����,�<� N�`�t���������̟ ޟ���&�8�L�\� n���������ȯܯ�}Ee�TM  [d�(�:�L�^�p��� ������ʿܿ� �� $�6�H�Z�l�~ϐϢϜ�d�SEV� ].�TYP�$��0�)߄m�1RSK�!O|�c�"FL 1Z�� ����߯�����0����	�:�TP5@����A]NGNA�M�$�E��k�UPSF PGI|%�1�%x��_LOAD0G �%Z%CAL�_TC� ���MA?XUALRM;'�@I(��~���#� V�#a��CQ[x�8��n���"�1060\	 �F�	�Ϣ������� ������ D'9 ze������ ��R=va �������� *//N/9/r/�/g/�/ �/�/�/�/?�/&?? J?\???�?k?�?�?�? �?�?�?�?"O4OOXO CO|O_OqO�O�O�O�O �O_�O0__T_7_I_ �_u_�_�_�_�_�_o��_,o��D_LDX�DISAc���M�EMO_AP]�E� ?��
  �5i�o�o�o�o�o�o��o��ISC 1]�� �oTd ��\no���� �����I�4�m� �f���$�������� �!��E�ƏT�f�:� ����ß�����z�� ܟA�,�e�w�^���� ��~������ �=� ��L�^�2��������� ߿�r� �Կ9�$�]��o�(t_MSTR �^�͂�SCD 1_xm�W���S��� ����=�(�:�s�^� �߂߻ߦ��������  �9�$�]�H��l�� �����������#�� G�2�W�}�h������� ��������
C. gR�v���� �	�-Q<u `r������ //'/M/8/q/\/�/��/�/�/�/s�MKC_FG `���/~��LTARM_2�a��2 ��#\`Y>G`METsPUT`�"�����NDSP_CMN�Ts506�5�� 	b���>�"1�?�4��5POSCF�7��>PRPM�?�8PSTOL 1c2}{4@p<#�
aA �!aEqOG]OO�O�O �O�O�O_�O�OA_#_ 5_w_Y_k_�_�_�_�_��Q�1SING_C�HK  +O$M/ODAQ73d
?�7�:eDEV 	���	MC:MlHOSIZEs0���eTASK %���%$123456�789 �o�egT�RIG 1e��� l��%��? �  A$�ÜfYP�a,u��cEM_�INF 1f>7� `)�AT&FV0E0�N�})�qE0V�1&A3&B1&�D2&S0&C1�S0=�})ATZ�� �H�E��q9m��xAu���X�������� ���� ��v�)���я��П �������*��N�� ���7�I�[�̯ן�� �9�&���\���� g�����i�ڿ������ ï4��XϏ�iώ�A� ��m�������߿�ѿ B����ϊߜ�O��� ���ߟߩ����>�%� b�t�'ߘ�K�]�o߁� ����(�_�L���p��+����������.ON�ITOR�0G ?�ak   	EOXEC1�#2345�`U789�# ��xxx*x 6xBxNxZxPfxrx22�U2�2�2�2�U2�2�2�2��33�3aR�_GRP_SV �1g�y�a(�Q���(?Y.���o�B���?��<l BHm�a�_Di�n�!PL_NAME !�5�
 �!Def�ault Per�sonality� (from FwD) �$RR2�� 1h)deX)�dh�
!�1X d �/d/v/�/�/�/�/�/ �/�/??*?<?N?`?�r?�?�?�?�?�?�82 S/�?O O2ODOVOhOzO�O�Ob<�?�O�O �O�O_"_4_F_X_j_�|_�_LhR� 1m�)9`\b0 ��_pb�Q @D7�  �Q?��S�Q�?`�QaAIڏEz  a@og;��	l�R	 0`4b@4c.a�P�Jd�Jd�Ki��K�J����J��J�4�J~��jEa�o�-a�@��o�l�@��z�b�f�@��S��a�Q�o�c��=�N��
������T;f��
���m��*�  �p  ��$p> p�$p��o?���?����{�����o�Bntr�Q�skse�}�l�p�  ��pu`j  #p��vks��� 	'� �� �I� ��  ���}:��È6�È=��9�N��b@^�d� �n�Q���{�R�x���nN. ��  '����a�`@a�@/�t�@p@p�nZ�CpC0�f0��+pB/pC3}�P��@%�Ea � oo$~|m����gAA%���. ���z�`�P���QDe���˟���(��m�� ��t O� �ru �4 ��R�c��s� �:�u�a�P�` �?�ffd�!���|��7� ��گ`쬛af��>搠���iP�P;�e�S�Ea<4f�u�>LX��s��b<	�I<g��<#�
<2���<D��<��a
vo��¯�S��S|.���?fff?u��?&찗d@T����?�`?U��?X����Z� ��T:z�TB��Wa�з *dů�ρϺϥ����� ���&�8�#�\�h�+�F. Kߘ�G߼�3����Wɯ���G�@ G����X�C� |�g�y��������� �jZ���ￏQ��� �ߙ�����3����� ��/A��t_�(��������� �d���@+FpA�IP�t��%���[`B�0�����<ze�cb!@�I�
�M`B@���@`�9@y��?�h�� �@�3�[�N��N�N�E?��<�/:/L ��>��ڟ�A��p�C�F@�S�b/DpX������@�t�?�%�h��`/q�G��Gkn�F&�Fצp�E,8{�/ F��ZG���F��nE�DE�,ڏ�/� ����G��F7��F��ED��.� �C?.?g?R?d?�?�? �?�?�?�?	O�?O?O *OcONO�OrO�O�O�O �O�O_�O)__M_8_ q_\_�_�_�_�_�_�_ �_o�_7o"o4omoXo �o|o�o�o�o�o�o �o3WB{f� �������� A�,�Q�w�b������� ���Ώ���=�(�@a�L���p�����(r!�3�ji��r���<ꕢ�3Ա�ڟ�y�4 ����y���P�2�D�&��jb^�p�1w���������ʯ����ܯ� �s�P^�PD�c�`�m���y�\������Ӱ�¿Կ� ����.�G���� }ϳϡ���홍�U�_�J���$�y.�@�v� d�z߈ߚ�x�4����@���� ��D�.�2� ;�$[�G�[�^��B���B��CH � ^����u�����������p�h�M�_��q����������"^�^�Y�m�2��
 ����#5 GYk}����p��h*�� ��>��x}��$MS�KCFMAP  ���� �����m�N"ON�REL  6��9_�"EXCFENBk
7]��FNC�}JOG_OVLIMkdu�yd"KEYk��"RUN���"SFSPD�TYU��v_SI�GNk}T1MO�T�z"_CE_GRP 1n��9\���/���/ �/4��/?�/2?�/'? h??�?C?�?�?y?�? �?�?O�?@ORO	OvO -OoO�OcO�O�O�O_��O*_<_#_`_-�"T�COM_CFG 1o/���_�_�_}
|Q_ARC_��6��UAP_C�PL�_�NOCH�ECK ?/ 5�;h9oKo]o oo�o�o�o�o�o�o�o��o#5GTNO_WAIT_LF'l5y"NT�Qp/z���q_ERR�!s2q/_�� R_���"�:�L�^dT_MO�sr�}, z�RP_��_�_PARAM�rs/������MW���� =e�345678901.�@�R� )�q���_�����˟��0��ݛLW�3�E��؏i�cUM_RSPACE,��������$ODRDSP��SI&�OFFSE?T_CARToݨ�DIS�ݢPEN_FILE�I!�Q��v�POPTION�_IO���PWO_RK t�'�C T�|�/�^�F�� ����Z���	 �m���A���i��_DSBL  Ķ�v���ޡRI_ENTTOj�sC���8=#�?��UT_SIM_D�J�6	��VàLCT u�}\���Q��W�_PEXE���RAT����� ���UP ve����������Ϭ*�8��$��2�#h�)deX)dh�>O�X dY�� �ߣߵ���������� !�3�E�W�i�{��� ����������2n�� )�;�M�_�q���������<����� +=Oas����X��� O��1m(?���(�.�g�}�"0 �д�u�  @D�  &�?��?р~H�D4  Ez�Z3;�	l	� 0ӀS@(SM� �i�i ��H)!H,��H8�Hm��G�	{G�8��6�MV��� �SC�)���)�����Ճ�*  �_p  � > ��  ��/$"��,��B,�Btr��«�H�¼	�/���/�"�#� �,0 �� ��  � ߽pj7   ��&X��?MU	'� �� 12I� ��  ���-=����U?g;/�@�}?�0~.ѱ�?;Ѳ����H[N �?A'�M�D�> C)�f)�" B& �"O4B+�<:�Q�@D1��oo$�_���JWAD0p�J@�A: �1 �E&?�O�O#__�G_2]�� ��t O� r�u �4 ���R�Uɳ� :�%Ёр� �?�ff��@[�_�_V_!{�o~��18р"oF0j>�P�Q6YPр�Zo�WrAdS�%��>Lw0�#�<	ƿI<g�<5�<�2��<D��<��׍�l�_��ѳMb�@?fff�?�0?&p:T@T��q?�`?Uȩ?X�-q �iyBq5Ya ��gI�_���� ��!��E�W�B�{� ��d�����ՏLnp�Ώ/�ʈG�@ G��U�ȏy�d����� ��ӟ�������yB =� ��?p���/򏸯 �߯R���'�9��o N�`�����~�����ۿ
ƿ�B�ĮD�e��ֿ;�ҿ_�J�?�A�h�oϨϓϸ��D4	��b!�_@���� �ħ��Ŀ����%�@I��)�M`B@���@`�9@y���?�h	� ��@�3�[N���N�N�E���<�/Y�kЖ�>��ڟ�A��p�C�F@��S���pX������@�t���%�h��߉!G���GknF�&�FצpE�,8{�� F���ZG���F��nE�DE,�ڏ��ૐ�G���F7��F?��ED��Mf�� b�M��q������ �����(��8�^�I� ��m������������� ��$H3lW� {������ 2VAS�w� �����/.// R/=/v/a/�/�/�/�/ �/�/�/??<?'?`? K?p?�?�?�?�?�?�? O�?&OO#O\OGO�O�kO�O�O�O�N(]�3g�ji�O�a��	U�E3Ա��O_<q�4 ��%_7_<q��P�Q_c_ERj�b}_�_1w������]�Y�_�_oP�_1ol��P�bPcn~���o�O�o{_�o�oY�`��o�o, /;M#�f0o�� ���Y�et�~�i#�1�C�yM�_����� ������{bS�Ԏ���	�?�-�c�Mj2����$�VG�z}�Bh����B��CH� }�9�֟�����0�B���wl�~��������Ư�T����\��qQ��U
 ί�0�B�T�f�x� ��������ҿ����܇��� ��]{x}���$PARA�M_MENU ?�Յ� � DEF�PULSE�	�WAITTMOU�Tl�RCV� �SHELL_�WRK.$CUR�_STYLj�Ϋ�OPT����PT�B����C��R_DECSNw�Te'�!� 3�E�n�i�{ߍ߶߱� ����������F�A��USE_PROG %P�%B��V�CCR��UeXÚ��_HOST !FP�!�����Tt`���������4���_TIME�� �T��  A�GDEB�UG��P�V�GINP_FLMSK]���TR����PGAʹ� |�[���CH�����TYPEM�Y�A�;�Qzu� �����
 )RM_q��� ����/*/%/7/ I/r/m//�/�/�/�/��/?��WORD �?	��	RS���CPNS�E̺�>2JO���BT�E���TRACEgCTL�PՅZ�� {`� ��a`{`�>q6DT� QxՅ�0�0}D�� #��Q�0���2%��Sc�0���2���2����2��2��2�4��4	�4�4�4��4�4�4 ��2��4�4�4�4��4�4�4�4(�4��2�4�4��
�2!�4"�4�?�?�? OO1OCOUOgOyO�O �O�O�O�O�O�O	__ -_?_Q_c_u_�_�_�_ �_�_�_�_oo)o;o Mo_oqo�o�o�o�o�o�o�m&�d' q 0BTfx��� �����7��%� 7�I�[�m�������� Ǐُ��1u�*�<� N�`�r���������̯ ޯ���&�8�J�\� n���������ȿڿ� ���"�4�F�X�j�|� �Ϡϲ���������� �0�B�T�f�xߊߜ� ������������,� >�P�b�t����� ��������(�:�L� ^�p������������� �� $6u�b t������� (:L^p� ������ // $/6/H/Z/l/~/�/�/ �/�/�/�/�/? ?2? D?V?h?z?�?�?�?�? �?�?�?
OO.O@ORO dOvO�O�O�O�O�O�O �O__*_<_N_`_r_ �_�_�_�_�_�_�_o o&o8oJo\ono�oV �o�o�o�o�o�o" 4FXj|��� ������0�B� T�f�x���������ҏ �����,�>�P�b� t���������Ο��� ��(�:�L�^�p��� ������ʯܯ� �� $�6�H�Z�l�~����� ��ƿؿ���� �2� D�V�h�zόϞϰ�������$PGTRA�CELEN  ���  ��������_UP y���љ������_�CFG z�)������<���� <�Z�l�<�$�D�EFSPD {�/��a�����I�N'�TRL |�/���8Lԃ�IPE_CONFI+�}}��Ѻ<�x�LID(�~�/��GRP 1���������@�
=�[����A?C�C
�X�C)��B��,r������dL�z��������� 	 �r�N��Ҩ�� ������B������������A���> ?�6>7�D_�������� ='�=)��������� 	B-��Q�M�<��  Dz����
��&L7 p[�������/�6/!/Z/���
V7.10be�ta1<�� B�=q�"`ff@}��">����!�=��͏!A>f�f�!@�ff�"��\)�"D��?��  �!@�!� �!A	p�#W��h/??*?�<?K;�w���� O/�?K/�?�?�?�?O �?O>O)ObOMO�OqO �O�O�O�O�O_�O(_ _L_7_p_[_m_�_�_ �_��_ o�_$oo!o ZoEo~oio�o�o�o�o �o�o�o DQy{/�#F@ {yw}� y{ջy�-����� �/�Z?l?~?w���t� ����я�������� �O�:�s�^������� ��ߟ�ܟ� �9�$� ]�H���l�~����_ۯ �����5� �2�k� V���z�����׿¿�� ���1�\n�j�|� ��������	�4� F�X�j�c�χߙ߄� �ߨ��������)�� &�_�J��n����� �������%��I�4� m�X�����ί������ ����!E0B{ f������ H�Zό�Vh�ϴ� ������ �2�D� V�O/�s/^/�/�/�/ �/�/�/�/? ?9?$? 6?o?Z?�?~?�?�?�? �?�?O�?5O OYODO }O�O���O�OtO�O�O _�O1__U_@_R_�_ v_�_�_�_�_�_"4 FxBo|����o ��o�o//0/B/; �__J�n��� ����%��I�4� F��j�����Ǐ��� ֏�!��E�0�i��O ^���N�ß՟����� ��A�,�e�P�b��� �������o o2oTo .�hozo�o�����o�� Ϳ�o
گ'�֯K� 6�o�Zϓ�~Ϸ��ϴ� �������5� �Y�D� Vߏ�z߳ߞ������� ���1��Uy�� :���������	��� -��Q�<�u�`�r��� ��������T� f�x�n������ ������7"[ Fj����� ��!//E/0/i/T/ f/�/�/�/�/�/�/? �//?A?l�e?w?&?�? �?�?�?�?�?�?OO =O(OaOLO�OpO�O�O ����*�O_@Rd�Z_l_��$PLI�D_KNOW_M�  ����A�TSV 킗�P�[?�_�_o�O&o�o#o\o�B��SM_?GRP 1��Z� �dI`�oo�$Cf�d����D��TPbj�o Lk�f�o"~�U�o> n2T�~�� ���7�4���p� D���R���ʏ������ ����6�
�T��*�������QMR�c��mT�EGQK? GR�� (�#���[��/�A�S� �����������$�� ��W��+�=�O����� ������� ���S��Ͻ�ST�a1 1Յ�����P0� @����E�ϲ� ��������M�0�B� T�fߧߊߜ������߀����7��,�m��2r�����A�<��z�3�������4 ���������5)�;�M�_���6x����������7����������8�(:L��MAD  ���� ���PARNUM  ���Ko���SCH�
 �
��S+UPD��xa�q{��_CMP_0�`� <Pz '�U��ER_CHK�����Z���RS8���_�Q_MO� ��%_��_RES+_G����� �� v/{/�/�/�/�/�/�/ �/*??N?A?r?e?w?J'��W,g/�?L%�� �?�?�?N#(��?OO N#w�4OSOXON#��sO �O�ON# �O�O�ON#�d �O__N"V 1�Uua�@cX���Pp�P$@cW���P��P@@cV���P�"THR_ICNR���pbA%d�VoMASS�_ Z�W�MN�_�SMON_�QUEUE ���e��`Ȩ`�N��U�N�V�2`E�ND4a6/NiEXE]oNeWBE\`>o/cOPTIO;g?+2`�PROGRAM %j%1`O_�~0bTASK_I���nOCFG ��o�9pDATA�ɓ�B{@ev2 w������z�� +�=�O��s����������nzINFOɓ��}�!dr��!�3�E� W�i�{�������ß՟ �����/�A�S�e�hw�҇ބ��| �9�8q�DIT ��Bׯj~WERFL�~hwS~�RGADJ� �ƪA�  �,�?E�8��Q�IOORITY�W���MPDSP�a�j�eU�WvT�OG���_TG���Rj��T�OE�P1�ƫ _(!AF�PE5 ����!tcp|��%�!ud�>?�!icm<�Q_n��XY_<q�Ƭ{�Oq)� *������Op������� �����<�#�5�r�Y� ��}ߺ��߳������z&�*�PORT�a��OpA%�_CARTREP~`|Ʈ��SKSTA�X^!*SSAV`�ƪ�	2500H8�09u�T毙䕣�*ƫ�����`X#��$�6�m�URGE�U`B��A)WFP�DO�V�2�W�q�?�Q�WRUP_DE?LAY �Ưe��R_HOT�hwR%�z����R_NOR�MAL�n��6S�EMI:y�Q�SKIP���X%�x 	����� ����X%-; %[mE��� ����!//E/W/ i///y/�/�/�/�/�/ �/?�/?A?S?e?+? �?w?�?�?�?�?�?O��?+O=OOO1U�$R�BTIF��NaRCgVTM�����m@�DCR�����ABnBzO��A�Q@��ާ������S{/ſ�8��?�*��æ���_]<	�I<�g�<#�
<2���<D��<��
+__{_�_)`�� �_�_�_�_�_ oo$o 6oHoZolo~oi_�o�o �o�o�o�o�o D V�_z����� ��
��.�@�R�= v�a����������� ׏�*�mN�`�r��� ������̟ޟ��� ��8�J�5�n�Y���}� ��ȯ�����A�"�4� F�X�j�|�������Ŀ ֿ�ӯ���0�B�-� f�Qϊ�m������� ����,�>�P�b�t� �ߘߪ߼ߧ������ ��(�:�%�^�A��� �ϸ������� ��$� 6�H�Z�l�~���{�� ���������� 2 Vh������ ��
.@R= O�s����� /�*/</`/r/�/ �/�/�/�/�/�/??�&?28�AGN_AT�C 1��K �AT&FV0�E02;ATD�P/6/9/2/�9p8ATA2>�,AT%G1�%B960k9W+++�?,�1H�?�,�AIO_TYPOE  EC/�4?REFPOS1� 1� K x	�O[H/O/�O �MNO`O�O�O�O_�O�C_�Og__d_�_+K2 1� KLON_�_�o�_*o�_5A3 1��_�_�_ o�o�o�o>@oS4 1�Woio�{o�o3W�oS5 1��o�oJ����jS6 1� ����]�H����S7 1��(�:��t��ݏ���S8 1�����Ϗ	���r����)�SMASK ;1� O  
���NɗXNO�?���1�.�8�1AMOTE � �.DN�_CFG� �U���5�0BP?L_RANGQ�K!�Y�POWER �Q5 a�SM_�DRYPRG �%�%R���ȥTA�RT ����U?ME_PROׯ��d�.D_EXEC_?ENB  �5]�GSPD=����Y3Θ�TDB����RM\ÿ��MT_ѐT���S�D0OBOT_NAME ��S�;9OB_OR�D_NUM ?���AH8�0�0I$�	���s	�\���ބ� ��e��	@̀}�D|��D0PC�_TIMEOUT��� xD0S232�n�1�Q; L�TEACH PENDAN��j�5���=Q�x0Ma�intenanc?e ConsK"-���"+�t4KCLS/C�}�6���|� No U�se�=[߹�F���N�PO�ќ�5�z_���CH_L@�3�U���	J��?MAVAIL`����+��]�I�SPAC�E1 2�=L ����p��扢�J@����8�?��� ���V�w� N�������������� �4�&G
l�}d	 Q5U1���������` 4&G
l}d(�#��2����� ���2A/b/%/ w/�//�/�3�� ��	/�/-/O/^??@B?�?�?�?�?�4�/ �/??&?�?J?l?{O��O_O�O�O�O�O�5 �?OO1OCO�OgO�O �_�_|_�_�_�_o�6_*_<_N_`_o�_ �_�o�o�o�o�o!�75oGoYoko}o+ �o�o����)��>��8Rdv�� H�����ӏ%�F�x-�[��G ��� R�;�
�� ����ԟ���
� �.�@����c���p���8�¯=�dؠ��ϟ ���!�3�E�W�i�_� q������x��կ� �'�9�K�]�oρ�w� �ϛ���Ͽѿ���� 5�G�Y�k�}ߏߡߗ���߻������ `S� @��8堯F�"�*ل����� �߇������,��� �V�h�2�<�N����� ��������.L 4v�R\n��Ĥ��
f�7�_M?ODE  ��M/S ���&�߂��Ïb��*	��&/�$CWORK�_AD]��x^�!R  ����t +/^ _INTV�AL]���hR_�OPTION�& �h�$SCAN_TIM\.�h��!R �(��30(�L8�����!��3���1�/@>.?���S22�411d�8�1�1"3��@���?�?�?���I-P���@����JO\OnOE@D� ��O�O�O�O�O�O_�_(_:_L_O���4X_�_�_��8�1>��;�o�� 1���pc]�t���Di�1��  � lS2��15 1 7oIo[omoo�o�o�o �o�o�o�o!3E Wi{����wc ���	��-�?�Q� c�u���������Ϗ� ���)�;�M�_�� �`[����ğ֟��� ��0�B�T�f�x��� ������ү�����$�7�  0��� o m��������ǿٿ� ���!�3�E�W�i�{� �ϟϱ�������v�� �/�A�S�e�w߉ߛ� �߿���������+� =�O�a�s������ ������ ��$�6�H� Z�l�~����������� ���� 2DVP�\�  �A���� ���%7I [m�����8��/ �/C (/N/`/r/�/�/�/�/ �/�/�/?F;/?�B?F�x1 �;?w=	1234�5678{�+�l�@�P�? �?�?�?�?O9/2O DOVOhOzO�O�O�O�O �O�O-/
__._@_R_ d_v_�_�_�_�_�_�O �_oo*o<oNo`oro �o�o�o�o�_�o�o &8J\n�� �o������"� 4�F�X�j�|������ ď֏�����0�B� T�f�����������ҟ �����,�>�m�b� t���������ί����(��6yI�[��@�`���������C�z  Bp*  � ���254F���$SCR_GRP� 1�(�e@(�l��0�@ `1 �[1s	 )�3�C� <�t�vrY�8P�}ϸkϤ����95C%����-u��ȡ����LR Ma�te 200iC� �190�1Շ0LR2C �3�=O���D�
f؜1u�2�U7��`1��v��@�u���	t����������$�^0� 2���_2T�gϡϊ�� o�F�D�f?��s������￶ht ,Z�-�r�B�˰�P�N��g�N�Aܰv�  @�DЎ�N�@����  ?� ��J�H˰��y��N�F@ F�` ������A,Q wb���n�N���������B� �_J�n�� ���/�%//I/ ��E+:3��6?|?�5�ա
�/�/�#��@=���"�/pǢ� 3Bm�07�590@7����EL_DEFAULT  I���� �^1MIPOWERFL  V�v5]2ރ0WFDOk6 �v5 �ERVENT? 1���O�t3�C�L!DUM�_EIP?�8�j�!AF_INExj0O�$!FT�?�=NOaO!Q�O ��PO�O!RP?C_MAIN�O�Hq��O�O�CVIS�O�I��OE_!TP&8PPU<_�9d4_�_�!
PMON_POROXY�_�6e�_��_XR�_�=f�_)o!�RDM_SRV�*o�9gouo!R�R8�o�4hdo�o!
��@M�_�<i�o!RLSYNC�4y8�oY!R3OS�?�|�4H� tO�8c����� ;��_�&���J���n� �����ȏڏ7�I���m�4���X����7I�CE_KL ?%��; (%SVCPRG1���안�!��3*�/��4�R�W��5z���6�����7ʯϯ�C�$�5�9��o G����o������ D����l��񑔯� 񑼯7���_��� ���4����]���� �������'��տO� ���w��%ϟ��M� ���u�������� ��?�A��Ͽ�ђ�؟ ꐊ���ɱ������� �?�*�c�N������� ����������) ;_J�n��� ���%I4 mX�|���� �/�3//W/i/T/ �/x/�/�/�/�/�/�/�?/??S?Ś_DE�V �9��MC:[8�i.m4OUT_Rf1~6~i8REC 1����f0�0 f0 �	 f0�2  
f0�4�1���3OMK�1�4=A%O^O�AA��
 �Z�6 s;B�3AA�qE=�=A���2WG�1*f0)f0{f0U�Of2}B0�����/Q�0�O_�5��@��@r�H�;@�  �x�0}@U@ܖ�O f0�f4�1aRf0�V_�2X0��@�f0?�@�~_�__���2\�0��0���0�@����_ �f0�f0�1=f0[Rf0�o�2T0��@�f0*�@u*oco�_ˌÆLH�0�0���R �  ѨRobmU�f0zf0娮o�2�Q��@�f06b�@z�ovo~K�LT=A�1(f0tf0�f0D�_c�f4e�=�ZZ� f0k0��0C�f0f0q��"~�N�LiI�1�2�f2P�f0>jI��zDf0bf0o.�g���φLU"f0i�0bf0��0���0V�b�f0jf0/f0|~ 0���E0��@�f0$��@Y�^�p���ՆL*��A�0=�Qpɀ�T�b�ʈ�f0_^�*f2C0��@��A01����&��2\�A4M��Up��A���p�<~��O��Ӧ�$X2�k�ҟ�2\&f0Z}��0�0Wf0��Z��b�f0f0RR~�[���F��@ݒq0"ޯ�*�a@� �Z�H�~�l������� ؿ������2� �V� D�zό�nϰϞ����� ������.��>�d�R� ��v߬ߚ�������� ��*��:�`�N��f� x����������&� 8��\�J�l�n����� ����������4" XFh�p��� ���0B$f T�x�����5V 1��<��FPs�\O�2 ѡ��A�5�a?_TY�PE�?k2HELL_CFG �z:f2/ HL�/<7RSա�/�/�/"? ?F?1?j?U?�?y?�? �?�?�?�?O�?0OBOVQK��p�!%QO O�O%��x�q�qQ��M��q�p�$�gBQ�d��O�O�&HK 1��+ �OE_@_R_ d_�_�_�_�_�_�_�_ �_oo*o<oeo`oro��oa&�#OMM �/�o�"FTOV�_ENM�t"!}*O�W_REG_UI��o�"IMWAITp�b���G${OUTv�$&yTIMu;��`VAL5's_UNIT�c�v})�MON_ALIA�S ?e�i ( he!� ��$� 6�%��c�u�����D� ��Ϗ�����)�;� M�_�q��������˟ ݟ����%�7��H� m������N�ǯٯ� �����3�E�W�i�{� &�����ÿտ習�� �/�A��e�wωϛ� ��X����������� =�O�a�s߅�0ߩ߻� ���ߊ����'�9�K� ��o�����b��� �����#���G�Y�k� }���:����������� 1CU y� ���l��	 -�Qcu�2� �����/)/;/ M/_/
/�/�/�/�/�/ v/�/??%?7?�/[? m??�?<?�?�?�?�? �?�?!O3OEOWOiOO �O�O�O�O�O�O�O_ _/_�O@_e_w_�_�_ F_�_�_�_�_o�_+o =oOoaosoo�o�o�o �o�o�o'9�o ]o���P�������s�$SM�ON_DEFPR�O ����:� �*SYSTEM*�  �l�*�R�ECALL ?}�:� ( �}6�xcopy fr�:\*.* vi�rt:\tmpb�ack��=>la�ptop-3jv�248ms:30�348 ��973� 3�̏ޏ�t}7z�a��������C�U���{�	�outpu�t\test_x�y.ls md:� over =>�3��0144:6�946�3�ğ֟�A{�����tp~���� ��;�M�_��6z����z����1�¯ԯg�?��z	�������L��^��9z�cal_dv����4�ſ׿�E����	�ʝ���L� ^�q�ϕ���4����� ���~� �2�C�U�h� zό�*߰��������π
�ߢ�?�Q�c���;�{�s:orderfil.dat�@���6������2��b:��遲����P� b�u�z�����6��� �������"���EW��8zߌԑ���3����C������ J\o��
���6� �����"��E/W/ j�|���2/�/�/�� ���/�/0��/G?Y?l��ptcp.pc@���6?�?�?�*5z?�0_1�?1�?COUO�?�?A2O#O5O�O�Ok?}?_�1��?�O I_[_� �1�V_ �Ef_�_�_�O�?_� �_DoVoiO{OO�_1o �o�ogoy�/���o GY��"/4� �j/|/?�/�C�U� �_�/��0�7�ȏڏ moo�o����A�S�e� �o
����џ�v �������O�a���� ��*�<�ͯ߯r����� ����K�]�p������ 8�ɿۿ� ���$����G�Y�f��$SNP�X_ASG 1��������� P 0 �'%R[1]�@1.1fϰ�?���%���Ͽ� ����� 6��@�l�Oߐ�s߅� �ߩ������� ��� V�9�`��o���� ���������@�#�5� v�Y������������� ��<`CU �y������ &	0\?�cu �����/�/ F/)/P/|/_/�/�/�/ �/�/�/?�/0??%? f?I?p?�??�?�?�? �?�? O,OOPO3OEO �OiO�O�O�O�O�O�O _�O _L_/_p_S_e_ �_�_�_�_�_ o�_�_ 6oo@oloOo�oso�o �o�o�o�o�o  V9`�o��� �����@�#�5� v�Y�������Џ��ŏ ���<��`�C�U� ��y���̟���ӟ� &�	�0�\�?���c�u� �������ϯ����F�)�P�|�_�x�PA�RAM ���}�� �	����P��p�OF�T_KB_CFG�  ����״PI�N_SIM  ��̶�/�A�ϰx��RVQSTP_DSB�̲}Ϻ����SR �	�� �& CAL_T�Cŵ�Ͻ�ԶT�OP_ON_ER�R  �����P_TN 	���A��RIN�G_PRM�� ���VDT_GRP� 1�����  	з��b�t߆ߘߪ� ���������+�(�:� L�^�p������� ���� ��$�6�H�Z� l�~������������� �� 2DV}z �������
 C@Rdv�� ����	///*/ </N/`/r/�/�/�/�/ �/�/�/??&?8?J? \?n?�?�?�?�?�?�? �?�?O"O4O[OXOjO |O�O�O�O�O�O�O�O !__0_B_T_f_x_�_ �_�_�_�_�_�_oo ,o>oPoboto�o�o�o �o�o�o�o(: Lsp�������� ��9�6�׳V�PRG_COUN�T�����d�ENB/�_�M��鴖�_UPD 1�	�8  
M����� ��-�(�:�L�u�p� ��������ʟܟ� � �$�M�H�Z�l����� ����ݯد���%� � 2�D�m�h�z������� ¿Կ����
��E�@� R�dύψϚϬ����� ������*�<�e�`� r߄߭ߨߺ��������\�YSDEBUG�n�Ӏ� �d��"�S�P_PASSn��B?4�LOG ��΅�� ����
�  ��� �
MC:\`��a�_MPCf�΅����ҁ��� ҁ��S_AV �i���l�� ���SV��TEM_TIMEw 1�΋ (J��F�����T1?SVGUNSɀo��'�����ASK_OPTIONn��΅������BCC�FG �΋O� 1H�2!`;A� I�r]o���� ���8J5n Y�}����� /�4//X/C/|/g/�/�/ ��,�/�/ ? ?�/�/H?3?l?W?�? ��?��0�?�?�?O �?&OOJO8OZO\OnO �O�O�O�O�O�O_�O  _F_4_j_X_�_|_�_ �_�_�_�_o�X�  o 2oPoboto�_�o�o�o �o�o�o�o:( ^L�p���� � ��$��H�6�X� ~�l�����Ə���؏ �����D�2�h�o�� ����ԟR����� .��R�d�v�D����� �����Я����<� *�`�N���r������� ޿̿��&��J�8� Z�\�nϤϒ���~��� ���"�4߲�X�F�h� ��|߲����ߤ����� ��B�0�R�T�f�� ������������� >�,�b�P���t����� ��������(��@ Rp����� ��$6ZH ~l������ � //D/2/h/V/x/ �/�/�/�/�/�/
?�/ ??.?d?R?�?>�? �?�?�?�?r?OO(O NO<OrO�O�OdO�O�O �O�O_�O__&_\_ J_�_n_�_�_�_�_�_ �_�_"ooFo4ojoXo zo|o�o�o�o�o�?  0BT�oxf� �������� >�,�b�P�r�t����� ����Ώ��(��8� ^�L���p�����ʟ�� ڟܟ�$��H��o`� r�������2�دƯ�����2��P��$T�BCSG_GRP� 2����  �P� 
? ?�  {��� w�����տ��ѿ����/�A�T�[��b�d�0 �p�?P�	� HBHA�L��|��@�B   C��`�϶ˀ��ϟ�D��F��A���x���A��qT$�9��6ff���f�@P�C�ώ�@�f߬��C��ߐ߮� �ޥ���%��%�D�W� "�4���j�|�����^��?Y�����	V3.00s��	lr2c��	*2�*�O�A� ��ї�33P�d��� qx�J�y�  �������T�JCFG [��l� o�V����������=K
%� Kq\����� ���7"[F j������ �!//E/0/i/T/f/ �/�/�/�/�/�/s��� ??(?�/[?F?k?�? |?�?�?�?�?�?O!O 3O�?WOBO{OfO�O�O P�<��O��O�O�O0_ _T_B_x_f_�_�_�_ �_�_�_�_oo>o,o NoPobo�o�o�o�o�o �o�o:(^L ������h� � �$��H�6�l�Z�|� ����Ə��֏؏� � �D�V�h�z�4����� ��ҟԟ��
�@� .�d�R���v������� �Я���*��:�<� N���r�����̿��� ޿ �&��>�P�b�� �πϢϤ϶������ ��4�F�X�j�(ߎ�|� �ߠ����������� B�0�f�T��x��� ���������,��P� >�t�b����������� ����&(:p ^����t��� ��6$ZH~l �������/ 2/ /V/D/z/�/�/�/ j/�/�/�/�/?.?? R?@?v?d?�?�?�?�? �?�?�?OO<O*O`O NOpO�O�O�O�O�O�O _�O__&_\_�t_ �_�_B_�_�_�_�_�_ "ooFo4ojo|o�o�o ^o�o�o�o�o�o0 B�oxf��� ������>�,� b�P���t��������� Ώ��(��L�:�\� ��p�����ʟ��� � �_�*��_�l�Z��� ~�����į�د� � 2���h�V���z��� ¿Կ濠�
����� .�d�Rψ�vϬϚ��� �������*��N�<� r�`߂߄ߖ��ߺ��� ����8�&�H�n�\� ���>�����x���� ��4�"�X�F�|�j��� ������������
 Tfx�D�� ����P >tb����� ��//:/(/^/L/ n/p/�/�/�/�/�/ ? �/$?6?��N?`?r?? �?�?�?�?�?�?�? O ODOVOhOzO8O�O�Op�O�O�O�N  P�S V$_R��$TBJOP_G�RP 2��E��  ?рW<RCS�J\��@0WP�R@�T�P � ��T��T �Q[R	 ߐBL  �UC�� D*W[Q�_�_�?fffe:l�B �P�ff@�`�33D  $a�U3o>g�_�_pox�l�P�e9<�bbY��?٪``$ol�oUA��gD�`�$�co�Quz9O�P�Aa�P@a���C�Z`Ep�o�]A6ffpu`aD9/�U�h�͔r� �~�a�RieAq�`�q�B�@9q�|�d&`8%���c333D�\P�8���?�`?L�pAp[QB�b�k�}�� ��z�� >�f9fԁL���T�f� �fo ��Nw@�*�8� f���r�,���П��ȟ ��'����F�`�J�X�X����SC�Vء���	V3.00��Slr2c�T�*��TQ�� �E���E�A� E��E���3E�iNE�!�hE�فEۑ��E�I�E���E���E�r�F�F��FM(F��5FBFa�OF�\F"�f,�z  E�@� E�� E�� E�  E���߫� E�����W EȆ�Ԏ�ᆰ�� F   F�� F$ F�j` F�@ F��P F�` 9�IR9�o����L�_ ���V��LQ�8TE?STPARS�X�UP9SHRk�ABL/E 1�J[4�S�V�+� �0�V�BV�V�WQV�	V�E
V�Vȥ�QV��V�V�뱅�RD	I��TQ�϶���������f�On߀ۊߜߐ�����ކ�Sl�RS  0ړ����������� �#�5�G�Y�k�}��� ����������/]k�o� ��*	�%�7�I������+�=�O؆�NUoM  �ETQ�PP �밆�_CFG �����Q@<PIMEBF_TTq��RS~��;VER�<Q�;R 1�J[
 �8�RP� �@5  ���� ��//&/8/J/\/ n/�/�/�/�/�/�/#? �/?Y?4?F?\?j?|?R{_�h@R
<PMI_CHANG� R �3DBGL�VQ`IR;Q�0E�THERAD ?U�E;@�S �?��?TO6V�0ROUT6e!JZ!�D�O~wLSNMASK0H|RSAA255.�E���O�O8TOOLO_FS_DIq��5�IORQCTRL� �s[���n]8 ]_�_�_�_�_�_�_�_ o"o4oFo�
�_Tofo��og�PE_DET�AIH3ZPON_�SVOFF)_�cP_MON �"�P2�iSTRTC_HK �J^mO��bVTCOMPA�T�h;C�d�`FPR�OG %JZ%CAL_TCP=<�n%QPLAYr��j_INST_M�@e �|�g�tUSe�]orLCK��{Q?UICKME�0)��orSCREF�>3Jtps��or �a�f��2w�_{����ZyISR_GRP� 1�JY ؛ 6���� �;�)�_�M��8�� ��Y�������͕�� ���/��S�A�w�e� ������ѯ��������=�+�M�s�	12345678�����f�X`�1�Ћ
� �}ipnl�/۰gen.htm�����0�B�X��Panel _setupF�}<��ϘϪϼ�����  u�k��*�<�N�`�r� �ϖ�ߺ�������� �ߝ�J�\�n��� ���I�?������"� 4�F���j�������� ������_�q�0B Tfx���� ���>�b�t����3�~U�ALRM�pG ?=J[
  �* /!/R/E/v/i/�/�/ �/�/�/�/�/??<?~�SEV  ��n6�ECFGG ��m�6��A�1�   Bȩt
 =?�s3E�?�?�?O O+O=OOOaOsO�O�G4z1ʂ��k SΟ��OH7Isv?}{�`(%0?"_p_I_4_m_ X_�_|_�_�_�_�_�_`o�_3o�L� �M��OAoI_E�HIS�T 1��i  �(�0 ��(�/SOFTPAR�T/GENLIN�K?curren�t=menupa�ge,148,2 Y,1}o�o�'{�+�o�eedi5t�bT��_Z�ouȇ�(.;M~CA?L_DV_X�o���*}-���sc�~�����)~'C��n7�1n�o� ��$�6��q,ǏU��pTCPn�@��������K��o8u����)�;�ʟܟ�a37��MV��������í�)a�a)o��� %�7�I�4sޯs����� ����Ϳ\����'� 9�K�ڿoρϓϥϷ� ��X�j����#�5�G� Y���}ߏߡ߳����� f�����1�C�U��� �ߋ���������Я 	��-�?�Q�c�u�x� �������������� );M_q �� �����%7 I[m��� ����!/3/E/W/ i/{/�//�/�/�/�/ �/?��/?A?S?e?w? �?�?�/�?�?�?�?O O�?=OOOaOsO�O�O &O�O�O�O�O__'_ �OK_]_o_�_�_�_4_ �_�_�_�_o#o�_Go Yoko}o�o�o�oBo�o �o�o1?�og y�����o�� 	��-�?��c�u��� ������L�^���� )�;�M�܏q������� ��˟Z����%�7� I�؟��������ǯ ٯh����!�3�E�W��Bz�$UI_PA�NEDATA 1��������  	�}�/frh/cg�tp/wided?ev.stmc����ҿ����)pri��.�Ip}2�V�h�0zόϞϰ� )���� �������0��T�;� xߊ�q߮ߕ���������Bv�� � *� �LT @�E�W�i�{����� ��6�������/�A� ��e�w�^��������� ������+O6 s�l�� ��� ������1C �g������ �L	///?/&/c/ u/\/�/�/�/�/�/�/ �/?�/;?M?���? �?�?�?�?�?0?Ot %O7OIO[OmOO�O�? �O�O�O�O�O_�O3_ _W_i_P_�_t_�_�_ �_�_Z?l?o/oAoSo eowo�_�o�o O�o�o �o+�oO6s �l������ �'�9� �]�D����_ o�oɏۏ����#� v�G��ok�}������� ş,�������C� U�<�y�`�������ӯ ����ޯ�-�����c� u�����������T� ��)�;�M�_�q�ؿ ��|ϹϠ�������� ��7�I�0�m�Tߑߣ� ����:�L����!�3� E�W��{�� ϱ��� �������r�/��S� e�L���p��������� �� =$a����}�r�����)�*��V hz����� ���.//R/9/v/ �/o/�/�/�/�/�/?��������$UI_�PANELINK� 1����  �  ���}1234567890_?q?�? �?�?�?�4��]?�?�? OO1OCO�?gOyO�O �O�O�OYIY0:�M���[0  SOF�TPART/GE�NA1?CONFI�G=SINGLE�&PRIM=mainedit �O�I_[_m_YJ_$_M=�wintpe,1 @_�_�_�_�]�_$o6o HoZolooo�o�o�o �o�o�o�o
2DV hz����� ���.�@�R�d�v� �� �����Џ���~�M 0,  9P E=Por?S�5�co:�{�^������� ͟ߟ��'�9�� ]�o�R����O�O���� �Z1�/�%�7�I�[� m�`C�������Ϳ߿ 񿀿�'�9�K�]�o� �L���э͙�S���� �������#ߒS;�M� _�q߃ߕߧ�6����� ����%��I�[�m� ���2��������� �!�3���W�i�{��� ����@������� /��Sew��� �.���|�# G*k}`��� ���/�1/C/֤ �͡�ۯ}����/�/�/ �/�/?�2?D?V?h? z?�??�?�?�?�?�? 
OO�ϝϯ�dOvO�O �O�O�OE�O�O__ *_<_N_�Or_�_�_�_ �_�_[_�_oo&o8o Jo�_no�o�o�o�o�o �oio�o"4FX �o|�����e ���0�B�T�f�� ��/���������ُ ���>�P�3�t���i� ����Ο��O/�s/(� �/L�^�p��������� �?ܯ� ��$�6�ů Z�l�~�������#O5O GO�� �2�D�V�h� ��Ϟϰ�������u� 
��.�@�R�d�v�� �߬߾������߃�� *�<�N�`�r���� �����������&�8� J�\�n���������� ������m�"4ßX jM�q���� ��BT7x ������A��/ /,/>/P/C�t/�/�/ �/�/�/�/o/??(? :?L?^?Ϳ߿�?�? �?�?�? OO�?6OHO ZOlO~O�OO�O�O�O �O�O_�O2_D_V_h_ z_�_�_-_�_�_�_�_ 
oo�_@oRodovo�o �o)o�o�o�o�o *�oN`r��� ��m��&�8� �\�n�Q���u���ȏ ������"���?�?��{��$UI_P�OSTYPE  ��5� �	k�{��_QU�ICKMEN  ���j�����RESTORE 1ו5�  ���/
�2�D�h�m c�������¯ԯw��� 
��.�@��d�v��� ����W���˿ݿO�� *�<�N�`�τϖϨ� �����ρ���&�8� J���W�i�{��϶��� �����ߡ�"�4�F�X� j���������� �����y�+�T�f�x� ����?��������� ��,>Pbt�� ����( �L^p���I���� //��SC�REܐ?��u1sc-�uU2M$3M$4M$5M$�6M$7M$8M!��UGSER/ 4/F"T. �O#ksW#�$4�$5*�$6�$7�$8�!���NDO_CFG �؜�  ,� ���PDATE ��)�Non�e V��SEUFRAME  
���&,1RTOL_�ABRT7?��N3E�NBX?I8GRP �1�!��Cz  A��3�1��?�?�?�?�?FO"OG:�ېUx81g;MSKG  {5�Ag;N41%a��B%��O���VISCAND_wMAXyEI�c8��@FAIL_IM)Gy@f���#�8�@�IMREGNUMryG
�KRSIZyC�,���$,SO�NTMOUW0{D��%�VU�#�c�� �P�2F�R:\�O � �MC:\XS\wLOG�VB@4 !�O�_�Q�_o
��z MCV��_�SUD10fE�X9k
�f�wV�2�ꜙ�p(��=��͓o��j�o�o�o �o�o�o�o 2D�Vhz��KPO6�4_?S�0��n6�uQ0LI Q�z�xr�qV� �|f@�w��� =	�xSZ�V�~����wWA�I��DSTAT ܛ;�@�_ď֏��$����EP12D�WP  ��P G/����q�AP-���B_JMPERRw 1ݜ�
  � �2345678901�������ʟ�� ϟ��$��H�;�l��_�q����LT@MLO�W���P�@�P_TI�_X�('�@MPH?ASE  53���CSHIFT�UB1~k
 < ���Ob��A�g���w� ��ֿ��������� T�+�=ϊ�a�s��ϗ� ���������>��'��t�K�!��#ޛ:	�VSFT1�sV:�@M�� �5��4� �0��UA�  �B8���Ќ�0p������Ҫ��e@��ME*�{D�'���q��W&%�!�M�$�~k���9@�$~�TDINENDcXdHz�AOx@[O��aZ��S�︕��yE����G ����2�������<���RELE�y?�w�^_pVz�_ACT�IV���H��0A ���K��B#&��R�D�p��
1YBOX� ��-�����2�D�1�90.0.� 83v��254��2�p�&���robo�t�ԟ   �pN g�pc� �{�v�xx���$%ZABC�3�=,{�낆;- !/^/E/W/i/{/�/�/ �/�/�/?�/6??/?$l?!ZAT����