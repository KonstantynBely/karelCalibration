��   ��A��*SYST�EM*��V7.7�0107 10�/3/2018 A   ���	�BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG,��DNSS* �8 7 ABLE�D? $IFAC�E_NUM? $�DBG_LEVE�L�OM_NAM�E !  ��ETH_FLTR~.  $��   �FTP_CTRL.� @� LOG_�8	CMO>$�DNLD_FIL�TE� � SUBD_IRCAP"� �HO��NT. �4� H�ZADDORTYP� A H� �NGTHph���z +LSP D� $ROBOTyIG cPEER�ބ MASKaMR�U~OMGDEV�l� RDM*N�DIS��� OTCPI�/ 3 �$ARPSIZ�oK_IPFpW�_MC-�F_I�N0FA~LAS�S�5HO_� I�NFO��TEL�� P�����R WORD  $ACCE� �LV�$TIM�EOUTuORT� �ICEUS��   �$O# ? ����!���
��
� VIRTUAL�/�!'0 �%_
���F��a�� 22+5�'�� =��!�!j?�����;  x?�5�=2~;#"oSHAR� 19  Pf?O(4OHO7OlO/O�OSO �OwO�O�O�O_�O2_ �OV__z_=_�_a_s_ �_�_�_�_o�_@oo ovo9o�o]o�o�o�o �o�o<�o`# �G�k���� �&��J��n�1�C� ��g�ȏ��쏯��ӏ �F�	�j�-���Q��� u����ן�ϟ0��7�z _LIST 1}�=x!1.k��09��j�1{���255.��r���	�05i�2p���砖�����̯ަ3诂�_� � �2�D�ަ4`���@װ��������ަ5ؿ���O����"�4�ަ6 Pς���vψϚϬ� c�$��Q>�$% =,8+5U�o!R�u�)��0H!� �����rj3_'tpd��31 � �!!KC� �߿�x(�'6��!C� �;�����!C�ON� ������s'mond���