��   �S�A��*SYST�EM*��V7.7�0107 10�/3/2018 A   ����SBR_T �  | 	$SVMTR_ID $ROBOT9�$GRP_N{UM<AXISQX6K 6NFF3 �_PARAMF	�$�  ,�$MD SPD_L�IT  �$$C�LASS  ������ � � VIRTUAL�\�'  1 �� � 8����LR Mate _200iC���BiSR1/�6000A���	H1 DSP1�-� ��	P02�.01,  �	���PaR�$ �� 8�w��M�������
=���r��r���9"�� � ����  ���� 2� E�r��  u��_ kk������ Q��!� 2{(���=���4 �= ���c	1�����&�  �5 ������ ��������� w��������2&�� ��9%�� 2� (U_!�N :?}q�� T`�/�/�/�/���/� ??%?7?I?��2��$���>��` �( �H 2�%�i0�-�� �_ ��>"�?�?�I%72A�zK]o�8E"{~;A�8r�����VT�{ $�����-�� � 1��4���?:��= � � [lq:��+�
= ��ʿ �$ͥ?5$_ =j?'5��M/_/ q/���/T_f_x_�_�/�_��3�_�_�_o����@�B> ���@U�FB}X'`X �o�Vo�4 "�?N�10.5�<=3A�J OO n ���_�K{n<D�� ���b
�	QG8CffH2e� ~&$��?u�3l��v��� � � `���r�[�M�� �����$x]o5$� ��?'��_  �c9	`R�%Q��x"�����"�4�F��_j� �_������ď֏���L���qo�e4/5�m4A�a�o�I@a �b�d��R�ab1�k����m0��	z�{�s��t� 9 �7~���E��� 	������$�<'�5# d������|���� �z¯ԯ���S��? @�R�d�v���������R��)��e2�31�h5A2F�����j�m�pq����h�.�.?Rz3	y �wݑ.g�� �������� �� ��� f������5$�����内�;��q��x"���(�r߄ߖߨ� �����9���&�8� J�\�n�����B��76!��?9��K� �`9H`g.�qσ���9�ȶ�Ϲς��� � q !�����	$���� ��[7"�݆Ss7�I�[�m�6HZ l�ߐ�ߴ����� 2[7p����=UqQ�Q[7v	v�a p�����	// -/?/Q/c/u/�/�/�/@�/�/�/�/?<�? 9?K?]?o?�?�?�?�? �?�?�?�3oaO� ��qO�O�O�O�O�O �O�O__%_7_I_[_ m__�_�_�_�_#?�_ �_o!o3oEoWoio{o �o�o�?-OO�oCOUO /ASew�� �������+� =�O�a�s��_������ ͏ߏ���'�9�K� ]��o��u��o۟ ����#�5�G�Y�k� }�������ůׯ��� ��1���U�g�y��� ������ӿ���	�� ����3ϭ���џ�ϫ� ����������)�;� M�_�q߃ߕߧ߹��� ����K��%�7�I�[� m�������#�U� G��k�}�E�W�i�{� �������������� /ASew�� �߭���+ =Oas���� �)�;�//'/9/K/ ]/o/�/�/�/�/�/�/ �/�/?#?5?G?Y?� }?�?�?�?�?�?�?�? OO1OCO��[O� ���O�O�O�O	__ -_?_Q_c_u_�_�_�_ �_�_�_�_oos?;o Mo_oqo�o�o�o�o�o �o�oKO}OoO8�O�O m������ ��!�3�E�W�i�{� ������ÏoՏ��� �/�A�S�e�w����� ��	ҟş?Qc+� =�O�a�s��������� ͯ߯���'�9�K� ]�o���ݏ����ɿۿ ����#�5�G�Y�k� �ٟ�����!����� ��1�C�U�g�yߋ� �߯���������	�� -�?c�u���� ����������sϥ� ��`����ϕ������� ����%7I[ m������ G��!3EWi{ �����1��� g�y���S/e/w/�/�/ �/�/�/�/�/??+? =?O?a?s?�?�?�? �?�?�?OO'O9OKO ]OoO�O�O//�O%/ 7/I/_#_5_G_Y_k_ }_�_�_�_�_�_�_�_ oo1oCoUogo�?�o �o�o�o�o�o�o	 -?�O�O�O��O�O ������)�;� M�_�q���������ˏ ݏ���oo%�I�[� m��������ǟٟ� ��Y"�����{� ������ïկ���� �/�A�S�e�w����� ����ѿ-�����+� =�O�a�sυϗϩϻ� 7�)���M�_�q�9�K� ]�o߁ߓߥ߷����� �����#�5�G�Y�k� }��뿳��������� ��1�C�U�g����� �ϰ�������	 -?Qcu��� ����); ��Mq����� ��//%/��J/=/ �������/�/�/�/�/ �/?!?3?E?W?i?{? �?�?�?�?�?�?�?U O/OAOSOeOwO�O�O �O�O�O�O_/Q/�Ou/ �/�/a_s_�_�_�_�_ �_�_�_oo'o9oKo ]ooo�o�o�o�oO�o �o�o#5GYk }��O__�3_E_ ��1�C�U�g�y��� ������ӏ���	�� -�?�Q�c��ou����� ��ϟ����)�;� M��r�e����˯ ݯ���%�7�I�[� m��������ǿٿ� ���!�}�E�W�i�{� �ϟϱ���������� ��y�#ߝ������ߛ� �߿���������+� =�O�a�s����� ����;���'�9�K� ]�o����������E� 7� [�m�5GYk }������� 1CUgy� ������	// -/?/Q/c/u/���/�/ +�/??)?;? M?_?q?�?�?�?�?�? �?�?OO%O7OIO� mOO�O�O�O�O�O�O �O_!_3_�/�/K_�/ �/�/�_�_�_�_�_o o/oAoSoeowo�o�o �o�o�o�o�ocO+ =Oas���� ��;_m___(��_�_ ]�o���������ɏۏ ����#�5�G�Y�k� }�������ş��� ��1�C�U�g�y��� ���¯��/�A�S�� -�?�Q�c�u������� ��Ͽ����)�;� M�_�q�͟�ϧϹ��� ������%�7�I�[� ׯɯs��������� ���!�3�E�W�i�{� ������������� �/���S�e�w����� ����������cߕ� ��P�߽߅��� ���'9K ]o������ 7��/#/5/G/Y/k/ }/�/�/�/�/!�/�/ Wi{C?U?g?y?�? �?�?�?�?�?�?	OO -O?OQOcOuO�O�O� �O�O�O�O__)_;_ M___q_�_�/�/�_? '?9?oo%o7oIo[o moo�o�o�o�o�o�o �o!3EW�O{ �������� �/��_�_�_x��_�_ ����я�����+� =�O�a�s��������� ͟ߟ��_�9�K� ]�o���������ɯۯ �I��������k� }�������ſ׿��� ��1�C�U�g�yϋ� �ϯ��������	�� -�?�Q�c�u߇ߙ߫� '����=�O�a�)�;� M�_�q������� ������%�7�I�[� m���ϣ��������� ��!3EW���� �ߠ������ /ASew�� �����//+/ ��=/a/s/�/�/�/�/ �/�/�/??q:?-? ����?�?�?�?�? �?�?O#O5OGOYOkO }O�O�O�O�O�O�OE/ __1_C_U_g_y_�_ �_�_�_�_O?A?�_e? w?�?Qocouo�o�o�o �o�o�o�o); M_q���_� ����%�7�I�[� m���_o�_ȏ#o5o ���!�3�E�W�i�{� ������ß՟���� �/�A�S��e����� ����ѯ�����+� =���b�U�Ϗ�󏻿 Ϳ߿���'�9�K� ]�oρϓϥϷ����� �����m�5�G�Y�k� }ߏߡ߳��������� w�i�����y�� �����������	�� -�?�Q�c�u������� ����+���); M_q����5� '��K�]�%7I[ m������ �/!/3/E/W/i/{/ ���/�/�/�/�/�/? ?/?A?S?e?��?}? �	�?�?OO+O =OOOaOsO�O�O�O�O �O�O�O__'_9_�/ ]_o_�_�_�_�_�_�_ �_�_o#o�?�?;o�? �?�?�o�o�o�o�o�o 1CUgy� ������S_� -�?�Q�c�u������� ��Ϗ+o]oOo�so�o M�_�q���������˟ ݟ���%�7�I�[� m���������ٯ� ���!�3�E�W�i�{� ��鏲����1�C�� �/�A�S�e�wωϛ� �Ͽ���������+� =�O�a߽��ߗߩ߻� ��������'�9�K� ǿ��c�ݿ������ �����#�5�G�Y�k� }��������������� {�CUgy� ������S�� w�@���u��� ����//)/;/ M/_/q/�/�/�/�/�/ '�/??%?7?I?[? m??�?�?�?�?�? GYk3OEOWOiO{O �O�O�O�O�O�O�O_ _/_A_S_e_w_�_�/ �_�_�_�_�_oo+o =oOoaoso�?�?�oO O)O�o'9K ]o������ ���#�5�G��_k� }�������ŏ׏��� ��{k