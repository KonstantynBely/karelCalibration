��   ��A��*SYST�EM*��V7.7�077 2/6�/2013 A�   ��	��BIN_CFG_�T   X 	�$ENTRIES�  $Q0FUP?NG1F1O�2F2OPz ?C�NETG  �D�NSS* 8 }7 ABLED? �$IFACE_�NUM? $DBG_LEVEL��OM_NAME �!� ETH_�FLTR.� �$�   ��FTP_CTR�L. @� LOsG_8	CMO>�$DNLD_F�ILTE� � SUBDIRCAP"m� HO��NT.� 4� H�ZA?DDRTYP� A =H� NGTHph���z +LSP� D $ROB�OTIG cPEEyR�� MASKa�MRU~OMGD�EVl���RDM:*�DIS�BOTCPI�/ 3 �$ARPSIZ�oK_IPFpW�_MC-�F_I�N0FA~LAS�S�5HO_� I�NFO��TEL�� P�����R WORD  $ACCE� �LV�$TIM�EOUTuORT� �ICEUS��  F�$O# ? ����!���
��
� VIRTUAL�/�!'0 �%_
���F��dF��04+5�'�� =��!�!j?�����;  x?�5�=2~;#"oSHAR� 19  Pf?O(4OHO7OlO/O�OSO �OwO�O�O�O_�O2_ �OV__z_=_�_a_s_ �_�_�_�_o�_@oo ovo9o�o]o�o�o�o �o�o<�o`# �G�k���� �&��J��n�1�C� ��g�ȏ��쏯��ӏ �F�	�j�-���Q��� u����ן�ϟ0��7�z _LIST 1}�=x!1.k��09��j�1{���255.��r���	�05i�2p���砖�����̯ަ3诂�_� � �2�D�ަ4`���@װ��������ަ5ؿ���O����"�4�ަ6 Pς���vψϚϬ� c�$��Q>�$%  =�/5+5U�o!R�u�)��0H!� �����rj3_'tpd��31 � �!!KC� �߿�x(�'6��!C� �;�����!C�ON� ������s'mond���