��   ��A��*SYST�EM*��V7.7�0107 10�/3/2018 A   ����DRYRUN�_T   � �$'ENB � $NUM_P�ORTA ESU�@$STATE� P TCOL_���PMPMCmGRP_MASKZ}E� OTIONN�LOG_INFO�NiAVcFLTR_EMPTYd $PROD__ �L �ESTOP_�DSBLAPOW�_RECOVAO�PR�&J_ � 4 $TY�PENFST_IcDX�$_ICI�  �MIX_�BG-� G_�NAMc %$M3ODc_USdk�IFY_TId �KMKR-  $LINc �  �_SI�Z�K� ?. � $USE_FLGA���i�SIMA�Q�zQB
'SCANz[AX'+IN'*I���_COUNrRO���3!_TMR_cVA�g�h >�i��'` ��p&p�!�+WAR��+�$$CL�ASS  �S���!��5��5� VIRTUz �/� �'/ 
55��������C8�0�!J5��5I1&;��?�?�?�?�? �?�?O!O3OEOWOiO�{O�O�O�Oc?+ W?�
501 a���O__  W1�J0�C O 1&; 4%�On_��G1W1\_�_�_�_�_ �_�_o�_1oCo"ogo FoXo�o|o�o�o�oW1@@S��&=^9J0��0 -rJ16t,��
1 >q�o`r���� �����&�8�?? �c>qW1j�|������� ď֏�����0�B��T��$?T�1&9 K������ ӟ���	��-�?�Q� c�u�J�������̯ޯ ���&�8�J�\�n� ��������ȿڿ��� �"�4�F�X�j�|ώ� �������������� 0�B�T�f�xߊߕϧ� ����������,�>� P�b�t���߼��� ������(�:�L�^� p���������������  $6HZl~ ���������  2DVhz�� �&V