��  ë�A��*SYST�EM*��V7.7�077 2/6�/2013 A�Q  �����ABSPOS_G�RP_T   � $PARA�M  ��  �ALRM_�RECOV1   $ALMO�ENB��]ON�iI M_IF1� D $ENA�BLE k LA�ST_^  d�U�K}MAX�� $LDEBU�G@  
GPCOUPLED1� $[PP_P�ROCES0 � �1��URE�Q1 � $�SOFT; T_I�D�TOTAL_�EQ� $,N�O/PS_SPI�_INDE��$�DX�SCREE�N_NAME {�SIGNj���&PK_F�I� 	$TH{KY�PANE7�  	$DUM�MY12� �3��4�GRG_S�TR1 � �$TIT�$I��1&�$�$T�$5&6&7&8&9'0''��%!'�%5'1?'1*I'1S'1]'2h"GSBN_CFG1 � 8 $CNV_JNT_* ��DATA_CM�NT�!$FLA�GSL*CHEC�K��AT_CE�LLSETUP � P� HOM�E_IO� %�:3MACROF2R�EPRO8�DRUeNCD�i2SMp5�H UTOBACK}U0 � �	�DEVIC#TI\h�$DFD��ST�0B 3$INTERVAL��DISP_UNI�T��0_DO�6E{RR�9FR_Fa��INGRES��!Y0Q_�3t4C�_WA�4�12HGX�_D�#	 d �$CARD_E�XIST�$FSSB_TYPi�� CHKBD_S�E�5AGN G�� $SLOT_�NUMZ�APRE�V��G �1_E�DIT1
 � Uh1G=H0S?@�f%$EPY�$OPc �0L�ETE_OKzBU�S�P_CRyA�$�4�FAZ0LACIwY1KR�@k �1�COMMENy@$DGV]QP� h���AL*OU�B? , $�1V$1AB0~ OL�U=R"2CAM_;1� x�f$A�TTR��@0AN�N�@�IMG_H�EIGHyAcWI7DTH�VTCYU��0F_ASPE�CyA$M@EX�P;$� Mf�C�FcD X $�GR� � S!1U`BfPNFLIC`~d
�UIREs3��AO}MqWITCH}cJX`N.0S_d�SG0� � 
$WARNM'@f��@� sLI? �aNST� �CORN��1FL{TR�eTRAT@0�T�`  $ACC�1"p '|�'r�ORIkP�C�kRT�q0_SF� *��CHGI1� [ Tz`u3I�PpTYVD�@*2 ��P�`� 1zB*HED�SJ* ��q2�vU3�v4�v5�v6�vU7�v8�v9���qO�$ <� so�o�h�s1�PO_MO�R. t 20Ev�NG�8`TBA� 5c���A�����]@�����ϋP�0Ѕ*��h�`
P�@�2� �,p�J,p_Rrrqo@b+�J/r/�J�JVq@�Cj��m�g��usp6�qP_}0OF� 2 w @� RO_�̿�WaIT8C��NOM_�0�1ەq3���cD �;���2�hP���mEXpG��0� F�p%r
$cTFx�JF�D3Ԑ�TO�3&@U=0�� ��H�24�T%1��E�� �e��f��f��0CPD�BG;a� k@$ƢPPU�3�f1):��A�AX 1�d�UN�$AI�3BU�FuF����! |��`��`PI�*�Pr�Mq�M~�����Fr�SIMQS@��G��QE���:��[MC{� �$}1�JB�`S�}1DEC�������ܴz� �ě0CHNS_E;MP�r$Gg�=��@_��q3
p1_FP󔞡TCh�@`�b���q0�c}�y�G�� V`�AԂ�!!���JR!0~ԂSEGFRA.p�v 7aR�T_LI9N�C��PVF������Y���Q���)B����( '���f�e�S���Q���.0�p�B��A����SCIZC�ћ�z�T���g������QRSINF3��p����?�������؉���Lot��G��*�CRC�eFCCC �`+���T�h��mh�Sb�A��h�*�f��:�DȬd�c��C��PTA�����w@�撀��EVT���jF��_��F��!N&�G�� X�������1i��! 1��,��hRGNP��"0qF���R}�D���2}�LEWN��Hc6����C�K�L�A�dCx :�L��ou2����A6N`Co�$LGp��B�1aP��s@�dWaA?@���~01R���dME%`�јd�_RAs3dA�ZC���z�OkqFC�RH`X`F�`��}��,�ADI; � 6b� ���`�p�`�5cn�S�@1�7a�AMIP���PY8CU�MңpU��iQU� $�P��C�CG1�������DBPXWO�����p$SKt��2� DBT �TRL�1 ��Q0T�i� �P�DJ�4L?AY_CAL�1R !'PL	3&@�0�ED�Q5'�Q5'̡&��DB��1!�W�;PR� 
�1� 0�1" �PA�$�q$�� ��L�)#�/�#mp�0$��/�$C�!%�/rq e�PEqr�&�/�rqic!REp�"'�H �O)@7"$LF3#$�#xBП W;���FO[ _D0m�RO(@���u���j���3RIGGE�R�6PA%S���E�TURN�2RcMR-_��TU�`?�u0�EWM����GN�P��zBLA��E��/$$P#�CP� "��&@�Qk�C5D�mpD�A#�p4\1i�FGO_AWAY�2�MO��fQg��DCS_(<�QIS ����c �C���A����B�t �Cn��A"�FW���D'NTV@��BVkQ��@���S˳W�sU�J&�xU�� ��SAFE��ZV_SV6bEXC�LUl�����ON�LA��SY��Q�tOyTBa��HI_V/>M�PPLY_�a��VRFY_#�q�B<d�_ )0��_+�Ip �TSG3�tp�b݀�0  AM���a*����0���Vi.b%fANNU�N� rLdIDp�U�2~S@�`mija�rj�f	�pOGI:�"+��$FOb��׀OT@w1 ?$DUMMY���d�[!�d١�& �E,o ` 8�HEx�s��b�SB$�SU7FFI�@ (��@�a5�g6�a���DMSW�E- 8�8�KEYI����T�MZ1^ӌq�1�vIN�����ir. D޵�HOST? ! �r���t[ �t٠�tYp��pEM>���$��S�BL��UL��/ A�|3����T50~�!0 � $9��ESAMP�ԕF��������I�0��$SUBe�Q�� ��C�:��G�SAV ��r���G�C� ˇ�P�nfP$80E��YwN_B�1 0�`DIad�@O���}�$]�R_I��� �ENC2_S�T � 2
ԇ J����L�q~S�`;����!3��M�I��1:�p�4  L�3�M��0��0K�4'a��AV�ER�q��}�M�DSP�v��PC�U����\ì�VALU�ŗHE� ��M�I�P@���OPP7  ��THS ���6�SH�F�F􁳠dL��0�T��SC�Q�d�:�ETo�5zrF?ULL_DUY�da��0��O�w�h�OT����0NOAUT5O�!6�p$�\֤��cl�
�C` ��C���`!�L��� 7H *��L���n�b���$ �0P�˴��ֲ��[!��@�a��Yq��dq��7���8��9��0����1���1��1��1Ⱥ1�պ1�1�1��2R
�2����2��2��U2Ⱥ2պ2�2�U2��3
�3��3�����3��3Ⱥ3պ3*�3�3��4
� ����SE�"8 < ��~��`�;I�����/��QFE�0�0� �9 ,��Q? z@^ ?�А��ER@#���A��z� :�`$TP�?$VARI�<�n��UP2�P; �pq�TD��S|�1`3�t���e�BAC�G< T�pr��)�p�bP�P o�IFI)� P ���U���P��P���0��� =t �;'�Ԡ��P'�ST (&�� &2&�r0E��*��	%�C��	��� _Cr�N�r��B��p�h�FORCEUP%b^n�FLUS�`H�N �E�h�RD_C�MK@E(����IN�_��&vPg�REMM�F~Q������ �3
K	N0�EcFF��N@IN�A��OVMl	OVA�l	TROV���DyT��mDTMX� ��m{@�
��? �*X[ ��CL��_:p�']@$�-	_
�;_QT��X
��@AQ	D� ��}��}!�V1� RQ��LI�MIT_�a椀�M���CLmd}�RIqV	�a��EAR��IO*PCC�����B�Bg�CM@��R{ �GCLF��G!DYM(/�aR#5TWDG��| s%�*�FSS& �s> P�a�!r1��EwP_�!�(�!1���E�3�!3�+5�&��GRA���?w�4�kPW��ONT��EBUG)S&2*�P|{@a�_E @:���S �TERM�B5AK5�`�ORI�G0BK6 �S�M_�Pr�G0CK6�U0A�9DK5��U}PB�E� -zA�a�@.PY3.@A$gSEG�:f ELEUwUSE�@NFI,��2�1ޠp4�4B�$UF6P�$�FQ4@�wAG0qTQ�&�HSNST �PATm�piBPTHJ�AߠE�p��2��P؀	E)�؁��1Rx�@�InaSHFT_���1oA�H_SHOR( ܣ�6 �0$�7�@9Dq�'�OVR#�naR�@I�@�U�b �Q�AYLO=�z��I�'"�oAj�!�j�ERV��:Qh��J��OG @@�B0����U����R!=P"�ASYM.�"�F�1WJG�уES��A�YvR�U�T @���E)�ᥳEP!�WP!��WOR @MB��G�RSMT�F�G1R��3laPA.@Q���`�q�uG � :����TOC�1�`yP�@ �$OP��ဝpՓá ��O,��RE�`RC�A�O�pтpBe�`R�mE u�h�A��e$P�WR�IM�ekRR�_�c4��qB H�2H���p_ADD�R��H_LENG�qByqnq�q�R��S.�I H��S���q�0Ӧu���u���u��S�E�'�LrS���J $��`��_OsFF��rPRM�� Z�HTT�P_�H�K (�^pOBJ?"ip��-$��LE`C!�Ƞ�L � �׬�AKB_~TS�s�S{`l��*�LVN�KR�n�eHIT��BG��LO�qt�fN�͂0���`���`SS{ ���HW��A�M�p�`INCPU�"VISIO�����+��t,��t,��� �IWOLN��N̠��C��$SLQb���PUT_�$��`{�P �V���F�_AS�"O��$AL��I����A��U�0��@Af��`q�<PH�Y���ÓZ���UO��#P `�����@�ڔ� �2�pP���`(�L��Y�B�Z�UeJ�Q�z�NEW�JOG-G��DIS�x�[�K-�f�#R �
�WAV�ǢCTR<�CǢFLAG�"[�;LG�dS ����Y�3LG_SIZ�o���������FD)�I�4�E�*�� D0���c$���𖶀����K���D0��� SCH_��߅p�2���N��F�T���E �"~�������U
�
�r{`L�	�DAU/ŃEA�-��dE�;�GqH�b�ᲐBOO��Uh Aɒ��I�T��y�[0ŖREC���SCR��ʑDeIēS.@��RGO� ��˒����d�´���	SU���W�Ĳ�Ľ��JGM$�MNCH|,�FNKEY%��KM�PRGK�UF�Y�PY�FWDY�H]L��STPY�VYذ@Y؀�Y�RS��H1`uۺ�CT���R��� �$�U	�m���
R��ݠғ`�G=��@P�Od�ڻŦ�M�F�OCUd�RGEX.��TUIK�I{�����	������I�M��@A�S�`���@������ANA���2�oVAILl�CL!~�UDCS_HI+4�`�s_�Oe�
!h�SȚ��|�S����IGAN4��F�J��T�bL� ��BUj � V 5!PT�$*��Hrv�Ϥ�e�@�AVrW !Pi�'��GP��1?2?3?�_� X � �i�=a�5���Ņ�ID$� tbP5R�bOh �Ĭ\A�ST	�RF�Y��0�@�  W$E�C�y����q_�� Y L� ؟0��@���`qFt�ǀ�FwҬ�_ Z �p����b��t�>0C��[ �p �CLDP	��UTRQLI{��T����FLG�� 1�O�1D�����LD���ORG�����췀hW>(�siT�r� 4\� �#0��վ�Sy`T�70y ' �$|�!�#RCLMC�$@B/T/�)Q��!=1I�p�_d] d�RQ>73$DSTB�p� c  6��-8AX�R� /8I<EXCE�S�b: 5Mp�1^��12�Td�2��0_�p"6_A:&��;�G?Y80K�d` \��GROU��t$�MB �LI9�CREQUIRDB�aL=O#KDEBUr� 1LYM��agbʑ`@p�C�"^MND���`c`b���̨�CDC���IN'��C��Z`���H��N�"�a#�� �EPST�� �c\rLOC�R!ITp��P�Ap��1 1ODAQ��d� X�ON�cF �R�fV�	X��b�U����u�1FX0IG}G�� e �y @X�a��X�XR�Q%��Y	��X	��V<�0ғDATA$`�E�a��a�N��f t $MDEaI:�)Sf��^d�![g�H5P�@]ez��a_cANSW�a^d�a��^eD�)BQz�� Xp�g �0CU4�V��`�=URR2{�h� D2�`A��A�! d$CALI&0ү�GS�w2K�RI�Nb�t<�NTEg�(i�bCu��=RBqg�_N�qjPukr����$ht�2kuyDIVF�&DHi0jp+�l �$Vp�C�$M�$Z�<!T �����b�emH ?�$BELT˪Z_ACCEL���;�"�IRCO�݁m���T���$PSi0�Lt�ڰW���Cp8��T�9�PAT!H���.���3]��Pl1_<�r��Ł�"S �Cr��_MG���$DD�9���$FW�`7`���.����DE�PPAB�Ne�ROTSPE!EՂ@L� JN�@�(0�t�$US�E_p�P&�ܦS�Y>��p�! �QYNr0A����OFFuan��MOU߁NGJ��܀OL~�ٔINC �d2Q��-2��� -2ENCSpa2U�X�+4R�IN�I]�0B����"n�VE��s>^�23_UPօp�/LOWL��[�` '���D>�2@Ep�]'��2C[pW�MOS���4MO��0�'PERCH  ��OV����蓼��� ���$�8S+�� 2@�������V�0^�O�L`�P��7O�U�UP"�8������TRK��AYLOA�J��1�����͵³3P� �RcTI�1	�� MO� O�-2�28 �`4�w�ٳ��?�pDUM�2��S_BCKLSH_C��P�ϐΦ ����bn�"�y�Ñ���CLAL V��!8��� ��CHK �SՐRTY����C��
*!6a_�ä_U�M����C���SC�L�W�LMT_J'1_L< 0-օa:�E4�U�G�D�J�P�J�SPCd�ȑZ���&3�PC �3�H_A@d���C� cXT��.�CN_rN���".�S��%�V���@:���ѹ�9���C' �SH�r�*�*! 9�9� p��^���9���3PA���_P��_�"�Ŷ�!ճ�����JG����~�OG|��,�TORQU��ON��޹*�B٢-�L*�L�_Wž�_�s�j��sj��sj�Ir�IJ��I�sFKP]�J�!X��c!�VC�0'42��1��{0��82���JRK��+� D�BL_SM���"Mζ@_DL�q�"GR�Vq�j�sj�sKH�_��I���
COS��LN- ��� ��p�	�p�	���ĺ�FZ� ٦KMY��D�TH�eT�HET0��NK2a3�s��s� CB�CB�sC&1n2���0��s��SB�s�N�GTS�1W�C.� 2Q�����$�'3$DU���8A!r �2P&�1Qb8V'$NE�4�PI� ��H�"%�v$�p�A��%�'���LPH�5�"h��"S��3� 33�"+3:2�pEV�(V�(�p�,V�*UV;V;V";V0;V>;VL9H�(�&�2P�-n�H;H;H";UH0;H>;HL9O�,�O�(O}I�.O�*O�;O;O";O0;O
>;O2F�"�Y��T�'SPBALA�NCE_T@SLE6�H_�SPHq��hR�hR3PFUL�ClX�R{W�R3Uz1=i
�UTO_�����T1T2�Y�2N ���`��Tq���Ps (d���T�O�p!�>L�INSEG����REVf��Q�DI�F��zy1j_g�r1k]�OBUa��t$y�MI`���SLCHgWAR>��AB��~u$MECH��Tˑ�a��AX˱P�y��f�'�r�Pl 
p�bI��:�ROB㠣CR��-u��ۊpM�SK_KP�tn P+ �P_��R��r_tn���18�c�a�_p�`�y�_p�aIN:a��MTCOM_C|���po  ݀�g`4�$NORE�S��r��`�rp �8U�GRJ��eSD�� ABג$XY�Z_DA�!F�r�D�EBU:a�q���pqu _P$��COD��G 1����`���$BUFIND�Xa�Hp"�MOR^Rsr $�qU&� ��u��ӑy�^��b�Gi�s � $SIMUL��8��x>���F�OBJEjP>��ADJUSψOAY_I��8�D����s�Ԑ_FIב=s�TZ��c�����`b�"�(�b`p0G�DN��FRIW�d�TgœRO%�A�Eb��HpOPWO> Vpt�0>�SYSBU<0[�$SOP��I�����U��b`PRUYN�rڕPArpDٖ��b��1�_OUT�Α�a�t$�IMKAG��\pv PDa3IM��1�IN[ �~0�RGOVRDY�˒���P�/�a�� �L_�PB�}����R)B�� ��MkᜪSEDb��` �N�@aM��~�Gq\�SLjP�Vpu x $OwVSLfSDI��DEX���q�����$o��Vb��N�A�@�'��,�'�D�M~y��]�_SETK�Vpv @U�^��ep�SRI��j�
q�_�}�����Hpdà*� w H\q�`���ATUS<�$T�RCx T�X�ѳBT�MڷıI��P�4p}Ѱ���Vpx D\p!E���β�0Ehbϱp�����ϱEXEհ@����)�=��f�ym��]p԰UP�L�$�`6�XNN����������� �PG�uzWUBñ�e���ñ��JMPWAI2[�P���LO7��p�FA`��$RCV?FAIL_Cwq�p��R9��p�c��(�}�x"�-�AR_PL���DBTB��,��pB3WD ��pUM*�"��IG�7��Qc�TNLW�"�}�Ry�iӻ��E�����Hp��DE�FSP` { L\p�`��_��Ճ�ӇUNI����Ѐ�RXD��Rb _LA`Pͱ]����pUq|-�#��q��O��XPc�N�PKSET�
��Pq��Uq} h�ARSIZE����=��u��S̀OR��FORgMAT�Pg�COנ,q�<bEM�d�����UX��,���PLI�b�Uq~  $>�pP_SWI�`���HqAXG�b�ALO_ o���A�r�B���C�rD���$EL���C_�lі� � � 1���r��J30 �r^��TIA4Z�5Z�6�rMOM��f���s���pB��AD`f��s����PU��NR����s��������Rt�� A$PI�&E�kqE�p- ~-�-�WC�0$��&�9q�gE���eSPEEDL@G �����Ծ����)� 9����)��	)���SAMWPx�0�1��MOVD�H$_S` Y%nk%_��1�t�2�t����c�v��8�H�PxIN��� ������(�+(+GAMM<Vu!�$GETE�U�ٓ�D5�
�PLIB�Rv���I�$HIBu�_L�ݰpB�&E�b�(A�.� �&LW�- �&�,�)	6�&1��f�`�j��� $PGDCK���ٓ_�����E���b7���a4��a9�� W$I��R�`D�c0�b~�Ե`LE�qkq0���81��0���`�Vp�P/aUR_�SCR��A�r��S_SAVE_D��,8Ex�NO5�C��y� 6�8@{$E�.{I��G	 {I�@�J�KP�q��H � ���x"Mao� ��s����d��6WP2U�Cqy���M� �k�F��aE�@�3�W<�@[�jQWg@���U�R�R��Sc22jQM"��[CL�W���M)ATr� � �$PY����$W`�fNG�O�`� b�b�b#�HЈ���a� ���c��X�O����Z�e��ހRt�# p䠰p�3+zO@�O�O�O�O�a5�_�r� |�E�8@��>v s�>v��8@_�kwVvy�AEހu%��"rB�\��P�"tP���PM�&�QU5 � =8*�QCOU�1 �wQTH#pHOL<�oQHYS��ESeF�qUE�p.BZ�O���  q�P���%��sUNְ�Q ��9OE��p� P2�3�p�AÔ�ROG�����Q2(�O}�2�������INFO�q�C #�e����RȾѻOI��� (�0SLEQ�с�рi�$C�{�D��L��`� QOK0r��!E� sNU!��AUTTA�COPYqu�?��`@ML�NI�M�X��Cᐛ� Y�RGA+DJ�q�i�X�Q��C$ഖ�`��W���P���0�������E-X8�YC0b�Ѫ�Obp�q���$�_NA9!��������`��� � Q���POR�A�.B�SRV0�)a�Y�DI��T_��{���@����������5���6��7��8y�*��PS8BL��m�M�C_F�p��PL9A8An�ȰR��9��р���$iB����d� ,�0FL-`L�C@SYN�[�M��C?��PWRc��L���!�DELA��8Y�5�AD�aAQSwKIP� �Q�Z4�OR`NT�� ��P_4��ַ@lb Yp������ ����Ƞ��ՠ���������9�1�J2Rܻ L�� 4*�EXs TQ%����(Q�����p�����p���RD�Cf� �`��X9�R�p�����r��~A$RGEAR_� sIOT�2FLG��vi��M%PC��B�U�M_����J2TH�2N'�� 1������G8 T00 I�����MlѺ`I�\8��REFr1�q� l�h��ENA9B{�(cTPE�0� 1���i�m���^QB#���:��"������2�ҙ����������
&�3�Қ7�I�[�m�(��&�4�қ�����������&�5�Ҝ�1�C�U�g�y���&�6�ҝ����������
&�7�Ҟ+=Oa(s�&�8�ҟ������&�SMS�K�q�|��a��E�?A����MOTEF����a@��L(Q�IOQ5�IcʦtR �W�0L�� �pZ����#p%�L���U�"$DSB_SIGN�1)Q%����Cl�(P1��RS2�32��b�iDE?VICEUS�,R>'RPARIT��D!_OPBIT`QY�OWCONTR;��(Q��O'RCU� M~DSUXTASKT3�N�p[0�$TATUn`P���RS�0RL����p_,PC9��$FREEFR�OMSp��%�GE�T�0�UPD(�A��2���SP� J���� !)$U�SA^���6���E�RIO�P@bpRY$�5:"_>@ �P}1�!N�6WRKI[D����6��aFRIENyDmQ�P$UFw����0TOOLFM�Y�t$LENG�TH_VTl�FI1R�`-C�RSEN ;IOUFINR]���RGI�1ӐAIT�I��4GXӱCI�FG2�7G1��Ѐ3�BƱGPR� A�O_0~ +0!�1REЀ�E3�e�TC���Q�A�V �G8��"J���u1~! ��J�8�%���%m��5�0G4�OX _0)�L|�T�3H6��8���%r4JE3GU�W�P�W�R�TD����T��а���Q�Tm�$V C2����1���91�8��02�;2/k3�;3 �:iva�9=i�aa��^S�jR$V��SBVB�EV'�V�BK�����&c�p��F�"{X�@�2q�PS�E���$.rRC��o$AŠFwPR��Gv]Ub�cS'�� 7�A6�I�� 0�@qV`��p�d`���E0�@���=�
B5S!� E��aRg����R��6�N AX�!$�A��0L(A���rTHI�C�1Y���h�t1T�FEI��q�uIF_CH�3�qI�G�a�pG1bxf���m����S@��_JF��P�R�ֱ�S��Ԁ��d �$SР��Z�GROU�̃TsOT�t̃DSP��JOG���#��_P��"O�����j��&7KEP(�IR���2�@M�R@�AP�Qn��E^�`�!�[�SYS�6��"[�PGu�BR�K�B �.��pIq��p��M���΂�`ADx�!̃9�BSOC׆��NӕDUMMY�14�p@SV�PD�E_OP�#SFS�PD_OVR=�b��C���OR�CNm0�F.����OV��SFR��pU���Fn��!#��C��A��"LCH����РOQV�s0��W�@M���ĥ:�RO�#ߑ�_��p�� @@�u@VsER�ps0OFSu@3CV? �2WD6���`2�ߑj2Y���TR�!����E_FDO>Y�MB_CM�D�B�BL�b>�f��attV"Q�240/p��N�Gg�z�AMx�Z�0���¿_M~��"7�<���8$CA�7�uD����HBK81,��IO�5���QPPA�=�"�M��5�͵���DVC_DBxC~� �3"�ТD�!��1��糖�3��@��pН�*��U�3��CAB��2VӠ�PѣIP��c�O��U�X�SUBCPU�r	�S�P P���90�^SQ׹c��."��$HW_C�Т��S���cA�A�pl$UN�IT��l��ATT�RI"���	�CYC=L��NECA��J��FLTR_2_F�I_�G(��9&�1LPx�?�>�_SCT�CF_��F_��6���FS8!����CHA��1�wᇲ�"v�RS�D�4"����q�_T��PRO��>�� KEMy_ܠ��8d��a d��a��D�Ib0!�RAILAiC��9RM��LOÐ C��Q*q��3q��V�PR��SQ�p�U�Cr�� 	�FUsNC��@rRIN'P`Ѹ0��u��!RA��B ����F�Ğ�gWAR~���BLQ�����A��������D�A����	����LD@)0��Q1�q��*q�1TI2rQǁ�p�$xPRIA1�"AFB�P�!|ߠ�p<`�R���MOI��A�DF_&@��51���LM��FA�@HR�DY�4ORG6 H����A�0 �MUL�SE&@"�Q��a ��G�	�����m$d$�1$1� ���0���� xm�EG�̃��`ARހ��09p�2o��z�AXE懗ROB�W�A��_�œSY�������S�WRI�@s1��STR�� ��:(�E�� 	%1����AB( �/&�a��ӰOT0^�	$ߠARY�sf"��ĚS@	�FI��*�$LINK���!%�a_%#�%{q�"XYZ82�*�qN�#OFF���"�"J�(j B�j�40С��n�3FI��%7`�q���j���_J�p��%��#�QOP_>$2H+5�3�PTB\12�2C��i�DU�&=62�TURN��2r��5t!}��p��|7FL��`���m�0�%+*7��	� 1�. K�M�&82�Q�2rQ�#�ORQ��G�� -(�+p��z�� 3q�E4"��T�GOV�@-A��M*�y�4�E:�E@�FW�J��G���D ��o�*� ��A7�P ��y��E�A�GZU:ZUL�CG�ER���	6�!E���B�TAFQ���)4����r'�AXУa2.q�c�W�c �W�c�W�p�Z�0�Z�0 �Z%@�ZK@�Z��Z
! �V� �Y� 
i� i�  *i� :i� Ji� Zi� �ji� zi�a�iDEBU{�$v�u��;q`��"F7O�50AB���6��CV�z� 
fr����ukњw�! �w�!�w�1�w�1�w%A �wKA�w��\0��".3LAB"2|Ew�x��҂�3 � E�ERVEN� w� $q�_NAǁ!_�PO����x` f�M�_MRA��_� d  T����ERR����~ T)Yi��RI�V"0�SN��TOQ�T)PL�H�T�ЅL�G�CJ_ � p�PTl X���_V1�b�Q���#�2�2+������/@��p��5�$W���V���VN�[�$�@�� �S���Q��	EHELL_C�FGN� 5�%�B_BAS��SqRvp0�K� �QS��Jϐ1a�%ΑU2�3�4�5�6�7�8�RaO���� � NL:Ɵ3ABn��АACKwv��)�o�u0�iႩ_PU2�CO,q��OU��P��ӕ`�����TP��_KAR�0��R�Em�� P����Q�UE٩��@���C�STOPI_AL zs��� �TĠ�� GSEM[�w�k�Mw�6y�TY��SO`��DI���Є�=�װ�_TMK�MANR�Qζ� E��$�KEYSWITCaH��Ѱ��HE��OBEAT���Ep�LE����&�U��F�d�����SO_HOuM� O��REF�@�PRi��R� ��Cr@�O0�p ECO��|�� _IOCM�4�M�k�K���'�O�# D�!ۧH�U��;��M7��@�3FOR�Cߣ�� ��O}Mq � @EtTxk�U#Po1B�TO�o3B�4x����NPX_AS���; 0ݐADD��(��$SIZߡ$�VAR�TIPRr�q�G�A(ҷ��@
�˨r�t�50�SV��XC����FRIF��R��S%�7�x���N�FѲEАO� x6�PSIڂTEC*�.%CSGL=�T�"�0�&�V�D��>�ST�MT
�o�P\�ByW�@?�SHOWw���P�SV� K�w� ���A00�0 �Q��K���O���_���Ti���5��6��7��8��9��A����@6������20��F�� 
 ����U ����� �����0�� �J@��:�1�G�1T�1a�1n�1�{�1��2��2��2���2��2��2�2��2 �2-�2:�2�G�2T�2a�2n�2�{�2��3��3��3���3��3��3�3��3 �3-�3:�3�G�3T�3a�3n�3�{�3��454��4���4��4��4�4��4 �4-�4:�4�G�4T�4a�4n�4�{�4��555��5���5��5��5�5��5 �5-�5:�5�G�5T�5a�5n�5�{�5��656��6���6��6��6�6��6 �6-�6:�6�G�6T�6a�6n�6�{�6��757��7���7��7��7�7��7 �7-�7:�7�G�7T�7a�7n�7�{�7��K�VP$�U�PD��  ��P���x�YSLO>��� � ��հ0�����QTAS�sTƠ��ALU}U�����CU��WFdQID�_Lѳ�UHI�ZI~�$FILE_Σ��T�$u�_VSA΁�� h��+`E_BLCK(�8bg�AhD_CPUQi��Qi����Sod_R1�ɢRw ��
PW,�d� �aLA�Sp���c�a�dRUN5� �a�d�a�d��5��a�d��a�d �T�pAC�C���X -$&qLEN~�3t���&p����Iѱ
�LO�W_AXI(�F1&q�T2mwM��ɢ�����I����Q�yT#OR.�&p�{DW��s�LACE���&p8�����_MAuйv8�u�w�qTCV�|��wTڱ�;�1�<ѷt���_��s��J����MD��ӠJ����u��
�u2q2�������l�s�pJKцVK~�hか��3ՃJ0����JJ�JJ��A�AL�����42�5Xr;�N1B�N�(�	��tL�p_k��x�"p��� `5`�GROU�PY�ӲB>$�NFLIC�ө�REQUIREv�EBUV�"q���кp2���#pɖ!qxг��� \��APP�RՐC���p
!�E�N�CLOz�,�SC_M ���A��u
!q޸�� 䣠MCp�r;�Xr|�_MG���C��,`��N��p��wBRK��NOL��t����Rϰ_LI��Hէ����JޠѤP� �p��p���p;��pD�"�p6�K��8��n�|"q���� Ғ�Mr:ql�Gqz�PATHv�������Rx��������pCNR�CaA��է���IN%r�UC�pwQ�Cd�U�M�Yop�����QE�:p�Gp�����PA�YLOAͧJ2L�HPR_ANqQ�L��`[�W�K�g���R_?F2LSHRё�LO\�䱕����ACRL_������޷C�XrH�P"�$yH���FLEX�� qJ%u� :2Dv�p4�K�GYq0�pPbt|F1Kљ� �׃�������E����/�A�S� e�w�����y���ф��@�蘏����J�ÊT���X����υ ��څ ��[����
�� �)���;�D�V�h�z�Y�J>��� � �������QIPAT��ё���EL4� �ؘJڿ��ߐJE��CTYRޱ��TN��F��ɗHAND_VB�p�ѹP`�� $�&�F2��K��ШRS�W9 qj��� '$$M��}�R��E@��Uw�H��sA�P H����Q���A���P
��A��Aɫ���j`���D��DɫP��G�`1)ST��9!��9!N̨DY�`���| �Y�鰋�KыǦ�J� ч�s�U�ХP�� &�/�8�A�J�S�=��� ; �t�.R66<N�/QASYM����	Ґ����Խ��ٿ_SH�����筈4@��+�=�O�JV���h�'CI����_V�I�dHN�u@V_�UNI�ÉD���J ҅�B�%�B�̦D�ųD �F�̓��������*U�c���Y��H̴`��XQENL� v�DIɠS�OwTqY�YP��� ��
�I�1A��äQ�`�Bc�S`�  p�a.a�o � ME����R'R�1TkPP�T�0) ���Qz�~� ��0�Xa	iT@�� $DUMM�Y1��$PS_f��RF��)$Pfm�aLA��YP��jb�S$GLB_T>mU�e�PpQ p���Q� X	�ɗ`��ST��ߐSBR���M21_V��8�$SV_ER��O�Ð�c�cCL�`�bA�5�O�RTPT O�P �� D �`OB���LO˰&uq�9c�`r�0�SYS�qADR�TP�PT�CHb � ,x&����W_NA��c�tz�9SR��?�l =�� M�u`�ys�u~�s ��s�������� ���0�)�T�"�5� ~���B����s�?�?�?|DY�XSCRE)�jp�ȐST[�Fs}�P!��t)�r _� Aq� T 	��`ob��a`�l��Ҩ���g�c�O� I�S�c��TX�UE��T� �ñjp^`S<q�RSM_iqmUUNEXCEPlV֑XPS_�a����޳�����޳R�COUx�ҒS� 1�d��UE�tҘR�b9�PoROGM� FL�o$CU�`PO?Q��д�I_�PH�� �� 8џ�_H�EP�����PRY ?��`Ab_�?d�Gb��OUS�� �� @�`v$B�UTT�RV`��C�OLUM��U3�S�ERVx��PAN�E� q��P@G�EU�<�F���q)�$HELPB�l2ETER��)_��m� Am���l���l�0l�00l�0Q�INf��SE@N0�� ǧ1��y��ޠ �)�;LNkr� ��`T�9_B���$H�b TEX�*��ja>�/RELV��DIP>��P�"�M�M3�?,@i�0ðN�jae���USRVIEWq�� <�`�PU�P�NFI� ��FOsCUP��PRI8 �m@`(Q��TRI}Pzqm�UNP��T� f0��mUW�ARNlU��SRT+OL�u���3��O�3ORN3�RA�U�6�TK�vw�V�I͑�U� =$V�PATH��V��CACH�LOG�נ�LIM�B���xxv��HOST�r�!�R��R<�OgBOT�s��IM�� gdS)} 2����a����a��VCPU_�AVAILeb��EX��!W1N��=�>f`1?e1?e1 n��S��; $BACKLAS��u�n���.p�  fPC�3�@$TOOL�t�$n�_JMPd� �ݽ��U$SSx�C6��SHIF ��S�P`V��tĐ�G�R+�P�OSURz�W�PRADI��P�_cb���|a�أQzr|�LU�A$�OUTPUT_BMc�J�IM���2��=@zr��TIL��SCOL��C����� ��Һ����������o�od5�?��Ȧ2ƢTEM�0�T9���vyDJU2Ѭ��� �WAITU��h��n���%��NE>u��YBO� �� $UPvtfa�SB�	TPE/�NEC��� �ؐ�`0�R6�(�Q��� $ش�SBL�TM[����q��9p���.p�O�P��MASf�_DUO�rdATZpD��J����Zp�DEL3AYng�JOذ� �q�3����v0��vx��,d9pY_���	��7"\��цrP? �QQZABC�u�� ��c"�ӛ�
,?  �$$C�������!N��P<� � VIRT���/΢ ABSf�u�1 ��%� ?< �!�/ �/??0?B?T?f?x? �?�?�?�?�?�?�?O O,O>OPObOtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo Zolo~o�o�o�o�o�o��o�o{� ��AXL�MT�s��#  �tIN&8qtGPREO��+vup�XuLARMRECOV �)Xrzu�jF �%�!d�� ����7�I�[�m�~�, 
�/��v�NG5� �+	 =#�
ڏ�� �PPLIC5�?��%upՁH�andlingT�ool -� 
�V7.70P/3�6 ��
]�_S�W2�D�F0j�W�� 43Y�J�9�K��7DA7?����
�&�X�e	-�NoKne��J�9p��~� �T7�	�_ ���_�Viu�6s��UTOz"�,tTy~.�HGAPON� �%��!.�U��D 1�y� t�x����y.�K�Q 1��{  Hp�������	���uq��"{�" �!���Hեw��HTTHKY��"ٯ ����u�����󿽿 Ͽ�����)�;�M� _�qσϕ��Ϲ����� ����%�7�I�[�m� ߑ��ߵ��������� �!�3�E�W�i�{�� ������������� /�A�S�e�w������� ��������+= Oas����� ��'9K] o������� �/#/5/G/Y/k/}/ �/�/�/�/�/�/�/? ?1?C?U?g?y?�?�? �?�?�?�?�?	OO-O ?OQOcOuO�O�O�O�O0�O�O���TOĀ���DO_CLEA�ND���{SNM  ɋ���_�_�_�_�o��_DSPDR3YR�_��HI!��]@�_}o�o�o�o�o�o �o�o1CU��MAX �bTQNQS��sqXbTB�o�B���PLUGGb�cWo��WPRC4`B�P]klo^�rO�r=o��/SEGF;�K�+� 6��_�_}�������ŏ�0�LAPZom�/� �+�=�O�a�s����������͟ߟ�6�TO�TAL�v�y6�USWENUZ�g� HX�L�NR��RG_STRING 13��
�M,�S��
��_ITE;M1��  n󝬯 ��Я�����*�<� N�`�r���������̿�޿��I/O SIGNAL���Tryout� Mode��I�npB�Simul�ated��Ou�tT�OVER�RW` = 100���In cyc�lHŕ�Prog� Abor^Õ�~>�Status���	Heartbe�at��MH F�aul����Aler�����'�9�K��]�o߁ߓߥ�  ^S��^Q�������� ,�>�P�b�t���� ����������(�:���WOR9���r��� L������������� *<N`r�������PO �������9K] o������� �/#/5/G/Y/k/}/�/DEV� - �/�/�/??)?;?M? _?q?�?�?�?�?�?�?��?OO%O7OPALT��^A��8O�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_�_�_LOGRIxp��a vO�_*o<oNo`oro�o �o�o�o�o�o�o�&8J\n�_*�R �ݦqo����� �(�:�L�^�p����� ����ʏ܏� ���PREGbNK��$� r���������̟ޟ� ��&�8�J�\�n���𒯤�����$AR�G_r�D ?	��������  	$��	[�]����.��SBN_C�ONFIG ���L�K�F�CI�I_SAVE  ��k�b��TC�ELLSETUP� ��%  O�ME_IO��%?MOV_H��¿�ȿREP�|��U�TOBACK���V�FRA;:\8� �8���'`��8�c�,�WINIa@8�^��,�MESSAG�z��������ODEC_D��}�C���O� ���,�PAUS!���� ((O ��J�\�F�|�jߠߎ� �߲���������B��0�f�t�%�*TSK�  5ݒϕ�/�UgPDT����d�����XSCRDCF�G 1��� �������&�8� J�\�n���\�n���� ������"��F�� j|����/e|�2�GROUN��|��UP_NAܰ���	2��_E�D��1
��
 ��%-BCKED�T-��}��p�g�Ӱ-2�p8��/�/�8���g2 ���E/��/��p/~/��ED3n/ &/�/J/\.�/"?�/�/ED4?�/?�/\.p[?�?5?G?ED5�? n?#O�?\.�?jO�?�?ED6ZOO�O6O\.p�O_}O�OED7�O �Ok_�O\.G_�_!_3_�ED8�_�o��]-�_Vo�_�_ED9Fo�_�o"o]-�o�oio{oCRoY_Vh��]1�{� LN�O_DELGE_UNUSE	�LAL_OUT� V��WD_ABOR���~��5�ITR_RTNz�ǀH�NONS)�������CAM_�PARAM 1�����
 8
S�ONY XC-5�6 234567w890Y �f��@���?�W�( А��8�h�хu�ڎ��HR5ǃ8��	��R570�B�Affފ����� �ڟ�ǟ�"���F� X�3�|���i���į!��CE_RIA_I�������F���;�Я ���G�P 1����s�����V�C���������CO�Ce ��(��ǀC8��e@��H��CCX��V��Ch��p��x��_�� C�����Ⱥ��+�=�G��ށ���HE/pONFI�G=�f�G_PRI 1�B�$r� ����������(�~�CHKPAUS��s 1���� ,wu j�|ߎߠ߲������� ����0�B�T�f�x�Њ���D�O����T��_MORG�RP 2?� �<\�� 	 �,� �P�>�t�b���5�����e�.�?a�a��D����K���d�P��V��a�- `�/A�

s��������b&�i\��ܦPDB������)
mc:cpmidbg���:�  -�-y����p�U   �  .s�/3� ��d�~��~��{C�Ve�/��/��{Qg�+/��/��{�f/s/i�u/�
DE�F �(K�)��b buf.tx�t�/�/��_MC*������d,53�����ʇ�Cz�  B�p�B���FB�8�B���~C� Cޢ��D3�u
q�D�zl'D:�"D�rBENNEA7EV�ߓ=�F�pgF=C��F�e,G����Gp��G�/��	ބ	6����S4����(D~������/��ʄ3@`à1zTB�D�V@�a  EI�5� F*� F�G�$ˀF[� G�R�kNGl��G���G��&H���G֓�H��߃]��  >�33 �ށN�  n^��@߂#5Y�Ed��A���=L��<#�
� ��_�*2R_SMOFS��.�^�9T1��DE 3��l 
 Q�;;�P  0_*_^>TEST�"__���R���#o^6C"@A�KY��Qo2$I��B�0�� �C�qeT�pFPROG %�S�o��gI�qRu����dK�EY_TBL  �6��y� �	
��� !"#�$%&'()*+�,-./01��:�;<=>?@AB�C� GHIJKL�MNOPQRST�UVWXYZ[\�]^_`abcd�efghijkl�mnopqrst�uvwxyz{|�}~����������������������������������������������������������������������������q���͓���������������������������������耇��������������������E��`LCK�l���`�`�STAT�c_A�UTO_DO���O�INDT_ENB;���R�QY�K�sT2����STO��~��TRL�`LE�TE�ފ_SCREEN j�kcsc 	��UπMMENU� 1i  <�l�ol�K�u� ��FS����柽�ϟ� ��R�)�;�a���q� ��Я�����ݯ�� N�%�7���[�m����� ��ɿ�ٿ�8��!� n�E�W�}϶ύϟ��� ����"����1�j�A� Sߠ�w߉��߭߿��� ����T�+�=��a� s����������� >��'�M���]�o��� ����������:�#p)+�_MAN�UALӏ��DBC�Ou�RIG�$�DBNUMLIM��,1e
�PXW�ORK 1k �_-<_N`r�wTB_�  m���Y0�_AWA�Y��1G�@b=�P�_AL� =��B�YҀ��`�_� � 1!�[ , 

:&d2/o/�&J�Mt�IZP�@P��#ONTIM�M�d��&�
�e�#MOTNEND��o$RECORD 1'kU2)?�!�O�?1-?&k�k? }?�?�?88�?�???�? c?O*O<O�?�?rO�? �OO�O�O�O�O�O_ �O8_�O\_n_�_�__ �_%_�_I_�_o"o4o �_Xo�_|o�_�o�o�o �oEo�oio�oBT fx�o��/� ����>�)�7�t� � pu�����-��͏ ۏ�����N�`�Ϗ�� o����)�;����� �8���\�˟ݟ���� ;�Q�گI���m��4��F�X��TOLEoRENC�B�	"��L�Ͱ CS_?CFG ( +x'dMC:\���L%04d.CS�VY�� cֿx#A V��CH�z� _/�x.�G��},��RC_OUT )��- z/��SGN �*��"��#��19-JUL�-25 13:0�8��27-wMAY��4:3���]� Z�t������x.����pa��m��PJP���k�VERSIO�N ��V�2.0.11~+E�FLOGIC 1�+� 	d���ٓ��p�PROG_ENB�2��WULS�' �p�_WRSTJN� ���"�EMO_O�PT_SL ?	��]�
 	Rg575x#?�74D�56E�7E�50i�dԂo�2E�d��j�"�TO  .����k�[V_� EX�d�%� �PATH A��A\��M�_��~+ICT�F��, '�`��eg��}�STBF_TTS�(�	��E��`���� MAU���ߧ"MSW��-D )��},t���.�!��]l�R�v������4SBL__FAULy�/�|�#GPMSK��^�"TDIA��0����`���!1�234567890xS�l�P��� ��//%/7/I/[/ m//�/�/�/�/�/LZ0PV �� �/�2?X?j?|? �?�?�?�?�?�?�?O�O0OBOTOfO8<x�U3MP$�I� �A�TR>�O�@PM�E���OY_TEM=P��È�3��4󜐰�DUNI	�w�Y�N_BRK 1���x�EMGDI_�STA	��_�LPN�C2_SCR 27[��_�_�_�_ �&�_�_o o2or�nSUQ13y_+?|o�o�oвolRTd47[�Q��o�o���_>P bt������ ���(�:�L�^�p� ������ ?Ǐُ�0� ,p��+�=�O�a�s� ��������͟ߟ�� �'�9�K�]�o����� ����ɯ�����#� 5�G�Y�k�}������� ſ׿�����1�C� U�g�yϋϝ�ׯ���� ����	��-�?�Q�c� u߇ߙ߽߫������� ��)�;�M�_�q�� �ϧ���������� %�7�I�[�m������ ����������!3 EW��{���� ���/AS ew������ �//+/=/wa/s/ �/�/�/�/�/�/�/? ?'?9?K?]?o?�?�? �?�?�?�?�?�?OK/ 5OGOYOkO}O�O�O�O �O�O�O�O__1_C_�U_g_y_�_�_�_�gE�TMODE 15v'Efa t�|�_GgRROR�_PROG %��Z%���HogTA�BLE  �[�1O�o�o�o�ZRRSEV_NUM �R  ��Q��`a_AUTO_?ENB  u�S�Zd_NO�a 6��[�Q�b  *U�6p�6p�6p�6p��`+5pOastH�IS�cYa�P{_A�LM 17�[ e���6|6`+t����&�8�J�x_\�bp  �[4q��R���PTCP_V_ER !�Z!6o�Z�$EXTLOGo_REQ�v�y��SIZ�܄TOoL  YaDz�r��=#�
ނ_BWDo�%��fQ���w_DI?� 8'E�t�TYa b[�S�TEPg�y��P��O/P_DO�v$v`�FEATURE �9'EQ��Q�Handlin�gTool � �DER En�glish Di�ctionary��7 (RA�A Vis"� M�aster����
TE0�nalo�g I/O��p�1
0�uto �Software Updateb�� "/�k�mati�c Backup~
�d
!���ground E�ditB�  25�LCame�raT�FX� "L�o��ellT��Lw, P��omm9��shۡ�h600���cou���uct���p�pane� �DIF���tyl�e selectvѡ- /�Con��~9�onitor���Hd�tr�Re�liabT�ϣ(R�-Diagn�os��Q�	�H�Du�al Check� Safety �UIFc�Enha�nced Rob� Serv��q ��v	ԸUse�r Fr���T_�i�xt. DI[O f�fi�� )��\�endܰEr�ru�L��  pr$נ*�rO�� @����ENFCTN_ Menuİv��.fd`�TP �In?�faco� � 
E�G��p;�k/ Excذg�C���High-Sp�eܰSki��  �Par+�H���m�munic��on�s��\ap��ur�f�?�X�t\h8yU���connZ��2Т !�Incr��str)�8���M-6�KARE�L Cmd. L���ua��}��B�R�un-Ti�En�v�(<�@�I�<�+���s��S/W�"�H�Licen3se���� ad����ogBook(S�y>�m)	���"�MACROs,~��/Offse\��f����H�!�Y�M�1�MechStop ProtZ��3� 5
�Mi�4�Shif\��B;6S�MixܰQ�����H�Mode �SwitchY�M�ok���.�� ��MTt�Q�g�� �5��?ulti-T����ܖ�)�Posj�Re�gi>���  ! ��PA�t Fun<1��6iB/��R��Num�Y�3�G�P�/��� Adju<��	�/2HS�)�� o(�8�tatu����AD ��RD�Mޱot�scove&� #e�v������uest 867.��o�\���?SNPX b��Y�<��)�Libr%�
�Ort I���� "����.S�o� ��s� in VCCM,����� j������㣀/I�� 7�10�TMILI�BX����g�Ac�c����C/2�T�PTX�� �Tel�n��Y@����K�P�CUnexc�eptܰmotn¾� ������\m725����w�|5���  h640SP CSXC��i � j*�� RI�N��We���50�,��vrl�زmcen" ��fiP-��a���P��Gri�d{�play F� O/��? ��EL�R;�|�20��O{RDK�sciiw�oload�41d�;st�Patd���CycT�h���or�iɰ:�7c DatMa� qu6�2�0��*�������FRL�amc�K�HMI De��(����k��PC�φ�Pass�word�644���Sp�����D#Y�ELLOW BO��	?1�Arc%�v�isu����#ti�O�p�^�! 2��a6O�po�� t��ֶcT1o�����HT���xy�	�  5 $�t۠ig��1�0Ơ 41\+�J�PN ARCPSOU PR+�8b!�OL0Sup�2fil� �!��E@-�;�7croc�82��v����$ 12jSS�0e4�tex-� �I�7�So��tf�ssag�� e��У�qP��,��� "Tc �Virt��v�!�����dpn�
�J�3�SHADf0M�OVE T�MO�S O TԠ�get_var ?fails l�>P�U~1E���� Hold Bus %��h��VIS UP�DATE IRTORCHMA A�|{�vYWELDTV �S ]�DtS: R�741��ouiPb�}�y��BACKG�ROUND ED�IT "RC$REP�TCD CAN �CRASH FR�VR 62z1�SC�ra��s 2-D���r ) "��$�FNO NOT {RE��RED �`� m ��JO� �QUICKaPOP� FLEN m4�1S�Loc��gRT�IMQ%�#�FPL�N: FG��pl �m�r`�MD DE�VICE ASS�ERT WIT gPCV;PB�AN#a�ACCESS Mo .pc��Jo���Qui±�Kbld�mgUSB$ ��t� & remov� Pg�SMB �NUL� ;a|�FI�X��C��ACHI�N,QOL�`MO �OPT ՠa��P�POST0�WDUs C�wQAdd�`�ad���0io�2֫�$P�`W\0.$�0`O�IN&�P:�fix CPMO�-046 isskueC�J/aO-�0n�r130Т- ���vRSET VAR?IABLES-P{�ޯR3D m��vi/ew d��M��&��ea���b��of� FD�5P:N@x� OS-1y0`�h� sc���t��s ft�lo��7 WA�P�Z�3 CNT0 1T�/"�ImR�)��ca �Pu��PO�T:Whenape=wB�STY E�{1�t��ptKQdo /GET_�p �p��VMGR LOl�REAd0C~QW�~1��(�l�s�gD�EC�TpLpING /IMPR�DR(p+P�B�PROGRAM��ERIPE:ST�ARTU� AIN�-;�ӠM/ASC�IIzPÂOF L�q�DPTTB: �N�pML$me hP���`:x�mo&��allW`!�ӤTo�rc�A�U�HC�i�LpԸth�`n�@ �ch��/GEA�!�t�ou͐�RCal���k�Sign`� �ND�ԗThresh123��`��09p� : MSG_P�+0er  �Q�=Aܠzeron���0 H85��RI�mA�n�2D��rc:�0I��OMEa`�p�ONaP5�  נS�REG:FF-Д� �]�'���KANJI*��n��J��c�0as�n d�!OA im�mc �INISI�TALIZATI����~1wem�����dr+� LB A|�UWqminim�rec[�c!�R���}m$�ro -1>��S�ܰir��@ұJ�*1pdETw�� 5`?��I�ow u��< s_e 1lc��YbPM���p�Q���R`vR�&�lu\�3�Re �0�4q�q1#���m9 <a�arn���~��Box fo���*PRWRI�PW�S���v�09 F�pu�p�de-rel2 d�p� j��`━�betwe��IN�D Q���igE osnap|�us��spo TME��7TPD#�DO�p#a�HANDL 1\�k�`vR��ȀD�n�y�S�v�Yoper�abil� �T*�:� H � l\p��V�q�b�R�< p�a*�c&2O�`FA,�.�-QV7. f.v��[GT�pi�s���� ɠtmLin�e-Remark� �� RM-�` �W�#SPATH S�A+PLOOS U�IFc�+5f fig��pGLA����Vrp�������U�0the�r�V� TracD���tW�\b�s7���d�t�� n�@ I ���3:���dK�=y��it k8�d�wPayR![2]��^�1: g��s���dow�XQ��0I�S�q�qEMCHK EXCE C����MF +�Xah>�� 35\k��)���QBt���'b�d��[�c���e �`xk�S�� BUGrt��cD$`PETpȵ��f�c4��0XP�ANSI��DIG���@OoPmetTC�CRG EN��C�EMENT�A M�̀K {�`H G?UNCHG �`� �EXT�P�2�bQS��93 wP8�x�O�RYLEAKq � H5gyq�PLC WRDN R �sO /u�QSPE=p��G*�V ��$��tn720\3pGR�I��A�rT�PM�C ETH��pSyU7p�`  j5/^n�PENS�PN,���*P ont�`B�ROW�`!sRMVo ADDz CN �qDC���PT3 �ALA2@ ���pS�VGN EARLqY�R��ŰH57�GaJLAYҀEk (@M�PPD�p:*@H�S I`P��OUCH8���V�F�q�comH�x ���ERROR� DE� nJ��RO�C�URS8pI��Nx4q�-158n7��RSR xP#aU�p���Rqy�T�F�z�;�pk��t�� �gՂ�B�SY �RUNN�  a|�`�BRKCT�!�RO�p3@ \ap�SТ�AXxP���h�8+ q��ISSU�r} sPX�PTSI��K1M10_�I�PSAFETY Ck�ECK[��Á ������<#X�� ��TWD2�@�@�I{NV��D ZOp�5X��t�DUA=Ly� "M6�0�J"rF#�E��dPd?NDEX F�,t*UF�"Pʀ��0sFRVO117� A�PT6�KtqF�ALPTP247�7D6_�P�!;HI�G� CC�t;SNPX� MM��tq�d~�Vq�q#�
"��>DETEC�Tq*@RRU�qA�P�5p�9 y�)<9���7T��Pds� k�	���!Q���� t\4A�;A0�o2 "Ke@" 8@�HI�qXF8@4@H�PRDC"�
�aMB8@�IXF�b���zOX@8@����a�G}E�B�Ccs�cr�J8@�Ndctrld.�A�NZE�A�5��Q��!�`�Df�8@�`m�878�Q-z;� ��� rm`�i
��PR̠78�@�RI8@0q�Q ( ~\Mp��0t��!{B8@�\tQ<OX�St0�32hB3nO�Vtp�A�@gLCF�L��� �Rplcf���J8@�WTamai�E8@mubov2_miTA�O�S8@�U`T[tT�AqPr67�4xSShape GGen��8@j�I�[R�`�@8@T����%qc (u8@��II�^��Q~C�a�[8@;Ynrsug0�4� � 4�C�tMr68@�r5hB5��zVnretsp e"r�Po�wng0bGCRE�Ka�ޠ��DAT�E�k�creat.�q�M��a�oksqgtpa�d1P��(�tput�Zj�{�������܆2�8@����Q����sl�o��� �hex�H�TB�8�ď�ke1yH�8@�pmZb�NbR�u7A+�nrgc8@ UQ�pp�bUZ�dp0a�j921xSpl.Collأcq�\A�b�RNq�UA� (J�8@ip�_�WA��_�Y���a7hB7�ͦt�p[� "TCLSx9oKb��clskyht[��s�pkckZd ���$�TQ���dA�r�x�710a- KA�REL Use {Sp�FCTN9��a�7l�0s0a�� ( ���a��~C8@��MI���c8hB8"   ��8@ v	��v	   �lmatea99�qM����E�mcc;lm5�CLM;�� ��j��E�et���aL1M	�h�yasp,���?mc_mot�B�N���8@H����Q��su�'��Q�ȕ�䅮���j�oi#�ߕ��A_l�og�Z���trc�B����ve�ϓ�v���QWX��6�find�erxSCente�r F1�lSw52a0��ha6rX� (<�cr,�Q�Ձfi�Q  �NH0�I�ۡ���A8@�uL��tq�a "F�NDRVϳ���et�guid�UID �C8@���������TA@�nuf;��P�����C�B��_z�Ӡo��qG������l���f�ndrTY��2䁴t�cp"�,qCP MtF�}38@517��6s38�E��gf6 ��(��K��Q��-�X�L�A�tm6�P�� ���Q���	�����tm�Ĵ�b8@aej��TAiex���aP�Aa�ذ�cpr�m�A��l�_vars��
��dwc7 `TS��/�6��ma7A�F�Group| s�k Exchan�gJ 8@�VMASK� H5�0H593� H0aH5@� 6V� 58�!9�!8\J�!4�!2���"(�/���;OMI� `@a0�hB0�ՁU4U1#SAK(x2�Q�0I�h�ӂ)�mq�bWzR�D�isplayIm�Q@vJ40�Q8aJ�!(P��;� 0a���0��� 40;�q�vl "DQVL�D쌞�qvBXa`�uG�Hq�OsC��avrdqq�O�xEsim�K�40sJst]��uDd X@TRgOyB�Bv40)��wA~���E�Easy� Normal Util(in��K�11 J553m�0b2v�Q(lV40xU�)��������k986#8Uϕ�|�rP "NOR��dw d.a}oKksu�O�W����OY�W`�j0�6�H� �menuuyP6�Mx�`wRX�R577V��90 �RJ989F}�49b\�`(�fity�����e��<?��Vsmh`��8@��C0�Sv�q�8����w�pn "MHMN<��ޣx�Ay`�o��3�u�`f�І�x�t ��tRzQ��LV��vP�#tm���|I�1{oPx" �2|���I�3I/B��odstǏًmnx����}ensu_�	L<���h!!��Rt~��huserp��0Ҹ�ʐcM�_l�xP�oe��рpoper�����xdetbo /�l>�x���Ps$p��`���OPydspw�eb͓��z'R��u�Rr101&S՟{tb�`2�Z4�30������`4�
�4�5���KQ�m[T��dUCalG40`�Q)p40}������9;��DA��? v	LATA�umpd�\bbk7968��68c�f�bl�41969y�9и|�D���bd� "�BBOXêM��s�ched����m�s�etuM:�����ff���40��n�41��8��40q�col��|��1�xc�ؘ���li ��X�0���j��&�8��4 <�ro5�TP �E�#��ryK412r��;�(T+Q �Rec'�ʈ1Iw��84�����Ak97�1��71�;���p?arecjo��Q�NS�[T���dXra{il| nagek��M ,QT2 *� !(�ĜR%<x�80P!bh��p��4���4�yDgl�paxrmr "XRM�g�l�brf{���n���kl��9turb�sp��㧑- �l0s15	�g�625C� Mh�+���)89��	+��B6��o�ҹ��x�7�q40�����pd "TSPDx�=��tsgl��l�:dQ���8Bc1t���K�vrE�a�ܮ�����  ��!���21��`( AAVM� �2�0 �@fd� TUP him� (J545� l)�`8 616� %�VCAM� ��CLIO] (�0:�5& � (F\ MSC ��Rt"PBsSTsYL�D!28 :2�\ NRE F2h S�CH6pDC�SU tpsh ORSR �r�D!04�SEI�OC& \fxh 542 LEX"� ESETn�8!H ���sh8 7H �OMASK�Ø"7>�.�OCO*`x�!0�3"6�!/400:66�$ G639.6[8LC�H!6OPLGR70=3
5MHCR��0�C� (! �06�A.�f8!54
��00D;SWb 588�180� �h!37 88 K(D�"02C24��N�27 q9�25���2-6�05��9�PRST bB/FRDMES�!zB��930 _ N�BA  6� HL�B 3 (~!SMވ@ Con� SPgVC �8!20z���TCP ara�m\TMIL� A��@PACET�PTX �@p T?ELN 96��2�9�%UECK��r� UFRM et��P!OR ORP I{PL%CSXC�0�j�1CVVF l� FQHTTP �stA")�I#� CG�HP8ZIGU�I�0�hPPGS oTool� H8�@�djZ��!@�h!6�3�%�@32Q\�31� B�h!96�%R6�51�Rs�!53 oTFAD�R41��8"1 ��oo�"9:��41775�"/@�P�VCTO�@�U�!�sh!80�%PRXyY�R�!770 �b~8 885 ol3P2� L� аdi� �`�ڳh LCP{Q� T'SS �b�26:���^�@CPE �HT@�VRC~�tQNLy ��@002 %�b	0dis� �`7� <��a\0�T�`1 ��`en�b4 6582�`)FU02Q0Π�o`p�Ptu�r4 d$r5N��RU0p@�nse�QJp1 A�PFI[ Jp3�g3}4�g40 al�xrE1t44w466� ts U0  7v��0O��r5�e�p7 �p "sw�a61d:��r4��r5 Qp!wGr`�$�p8R�"s�P`tQ�b�36w717�w8`�v83���r�8�&:��pOq8�8 _"rkey8�9F�v�a90�91 p�p#@��� �D095�g[97*pur�A1@ d���P|P�q1�0QplSq1p#4��]a!sM1@sl༂8��H��\1�d1�`��v��@{�14p�ae��5# h2��`�6ޣ��7�f1p@��d�YpCq(d�ـd�1�`uq���� Cu1< Oq� ��7&ReU1$ �u1�Pϱ�� ��@- WQ1�58 ase C渒9 B��60 �82ń�p���4 (Wai��`吢!���7E��8�EU1&P`ro9�<�1��<�2��<�	0��T��"l�5J�l��cC���9%�MCR��P��2�`�Q2@96I7�Q��8��9Z�A2TPB���P�2P7�U5@�o���
�58�`U���3 w����?A�E�1��c�qAw�l��A�1��512# f��1�u5Р��"�a5p$��56�+aĈ�Q5h��Ұ�1 �@��pp�b[�538 xaB��|p�4Ⱅ2�11/q5�p�4U=5�P16 (߲�P z��0��8�P��H���p�e5`�e5(�/�P`bbf>�X��$�Z�U�5d�\�� X�7 	  ~��8 k_kv���79 s�82 &�H5��E6���p�����h���ñ���3�J"�`��4 3Ȥ5�9ѧ6�0t���8Ⲗ6D0$�$�4 7���!���<�j67?0\tchk<�P`s��<�B<�90���7�<���<�\K�<�q �Ӻ�A�C<���q�<д��<�t��sg<�lIc���FA<�H���<���<Я���<�hk ��<Щ�B<е�o�<����<��K�<�dflar��<Ш��� ��@o�`���D�;�<�gEvam����B<гoќ���<а�KЀ�creexl����P�`��<���|���j6<�=s��prs.`��� \���<�7������fsgn��P�b�t�at��<�L��1|B !�svsch/ � �Servo S΋�ule>�SVS��44�1u�_<���� (����ched��,��~��A\�� �� B���B�qA�h���cj�� � 5�1<���Ә�p��css "ACS <�&(��6� ������c el���Q�����torchm�s�<�- T�Ma�`Ѵ���09 J5�;598 J681s�7� 8��b���<Чa����te,s�����/�E��� m��ARC..�� 1q�4�!=�,�C�tc�pA�@t����f� F����7#�2x�SE�r����UtmS�09610'���RC�������� p��96`G= '��"H5W�@���L���\f� � �PATb���`!a4U�#!Stmt��E ��� �pM�A�!p��z�2?�i�n_<�X��r�X e/cW����V����etdl�vߏ\oveto���܏���mmonitr`�\��|#�0st��?.6a��PP�����! Q�!y`�`asme �Arol�6c�43�0 �pl���01� 25��  �<� v	�v	�A>@�818\n; <�s�I�B�2�pMPT�P"��C�1mocol��,��CT�v�'!`� �A���8P53��y`Touchs�s0�`��<��J5��@�Ѩ`mP����n[P Q�a,�E�a��IPL&
�Pth�A<�KF#xR�m;�Qetth�THSR'�q-�Rt���o "PGIO��#!$s�ISwka�"cWK��!�MHqWH54��5w5n/"�Sm/��@ 7�*�da��8`!w/Ac��tsnf Tk�/�#@gb�a��u`��^m�`Au��Zӭ�ܱQp��@��#���Ka<��M��t5QtZ�a<��d�FS5GK����G�1o1r��dW��64��tP@x���P ����x,� �?$���P<�Z4e�7�g "SVGN�.ox�copy "CO;�Wj$�O�A�9� "FSG�ѧ�%�7��_��f� wQS�WF*!"(�sgat�uɀ���_
��tpN_TPDo��9�79�#dߎ?���h��GAT���!#��  �Гf�` �@�"/� �w�Z� �b?6 ?� ����� ���E �8��M� �chrT� �K6K� �sms� �o6��ѐ�gtdmen�?3 �?��� ���mkpdtd2 ���, ���pdQ�X� ������ ���mvbkup�. �[�C�С��mk3uno��prp���Gmkl �4��s ��niU��� �ldv9rw���glg�4��� ��棑��aut7�.pб�旐 �ַ������su3� ��@�� �Ƿ� ���\ �6�b2X� ��&�� �x����A4�  ���B   946�" ��fB� �t\p�aic\p4k947 ���F#���� ��ictas���pa`���cc:�<��8o�����gen�� �I ��F�lnp � �Ď��stf@��1��wbO�c��Ջ�`��߄�vri�ߢ�а�-T� ���p�flo�w� OPAc��ow���R50qtS �#T� (A��4�#�0��pѣV�cu3�Q0F� ��SI�ac�����46����s&��p�a��!!���� ���55�b �o)�p���0�|��
�afcal3�P� ��f��}���`�f��m	߳�p�d�m�/���a/��$C`ѷ��� �! trac�k\P� 0�ine/Rail Tr��]TJ�69W�T  (L��8(`љT.�`� %��D��P0� (��8�48��_ɛ�₇�4����� �3b�b3���alV@ �NTf���%��I�in]0m���aen������&?5�8c@Itst3@�� $����`�,R9�%����0氱%��po�peners-OW dDev��F�M�6W���|A�Pc"�l!esv� �,��R�V$�Q���U<�V$ �k)9j �6��# ��ȼ��%paop/!O�PNU�V ��2c#elL��8g_��8/�6��tscG��$Ѐ�V!�3� 5vrCop�ߡ�7`�n( `�V"2D�a V'O$�:S9��� Pump E��jQ�@�" ��!
��@бMSC#�@��)P���AC�`��� � �v���� \mh/plug�@g�"�7P��uK")㠱io�7�CJ0��E�LI�O q1g 7A93շ�5 q9 t����]4rb ST��R�ÞCPJ989�P�L�SE�' �e C3Q(P �/Ov���o�P� ? I1�R����55��f�I1`�tcwmio��MIO������Utco1"CL�01V �cBK`iEo��uM?���Sl� I0�ߢ�Eg �o���fb �tI4\onfdtI����e%�p27�Inste�TB CoMIoo1E�R�(do554 (;r>Ex�,��nR##ipc��/>��qp5���
@oQé�1�p����7/o����ra�pd�CD V_��rP�֮��qp2Gcnd��s �p��a�o�r`҄�S��"�bc�a�c���2kI�<�?A�pcrt���or0�qd#��"���3p�+���D��Џ��vr2k�0���AG�.�+��cho�;�u�C��(� �uV630 �fwe P�mී�@�X��`��TX�� ��>d�chp "_��(	�3�����8����\p3�v�������9�3�1 ������low�[ͧ���c!hk���㳦s��s?Ө0�i�1h���2�� i�w����s?1*�`-	�:�O��vr�������0�'���PFR�APWat?1rn�eE�P�sp�& ac5�� _A�rbo#�, �a��g�������z�Qs<�ICSP+� 9_����� ��F�A9PH51�IQ93 7��HX6�hQ]PVR`S5��fPR�6 iQWPR� (�P!am S�u�"�A�I0�tppr�g�0���`h�@2atk932�!��E��^��asc "8�C8��S>i�atp�"��d�@1I�
g�ds�blfltJA�Qs�able Fau�P{C!��EV0ex~/!DSB (DC��t�$�p��X 7�@� �� 5��Q�t3*��~���td9� "`!%�(5��sb9������\	�6#���@�5�p$D@550-A�djust Po'intO"tVJ�Rs�z�䐄��!�X_�Yj���0\sg��4x��}7y�\ada�O"ADJ���j�Q�etsha<�SH�AP�sŭ'jpo �r4�t�!��$ �(�C|�	Tk!bRP�KAR/Qiagn/ostì!O!vV66 J`ew0��(�L���/�&krlde� ��PP�� �hU b���r3�Pyp?q��DBG2C��� �X�o�1U��� ��WT`�@i�pJCM�aipper Opv`1Se}�78 (MH G F� ;":�&##�� a��x�֕$��388�C�����#��9.�9�C��g##PPk�Q��8 �!�_"$�"��=0%�P� �A $��_�#%0AQ�C�~2 Mat.HandlE��!= &�pq MPLGET�0�1(�3�Tt&P�Sٰ' �B�1��B0����&p� �H��PP �'p��@�C 7PP	�TG�tD5�}�m�q�Afhnd �"F_R  ������PP	   pxT?Q���P(Pa���To�����?�p�mpaO��JP ak925��2`@O�JR	psQ`B2�unLHP�T7gse�GSo1�O�W�QT��v !�R��Ptp~���JRdm�on.�@��V�!ns�hYvr�QJ�g�Q`�o�jY�HS~7sl�f] ��pen�PDnRp(R&���ɐ823'� �ٔq���g� ����� 1�� S�� ? �c\sltQ�!|QE�P��a �rtPg��P�� �v��"SEDG8�s0.�qtdgY T�� ��vP`ho�s`<` ����qc�`g
�e`� o�w�a@o"�ile6�H�e�ȅnR��� �e! j517�>Ճ��J%��e�`��Q4��Q&�!L�!F�J�=�o�5�z/l17���_�œ���`C0C�  ���LA/NG j��A��p������gad����#�jp�.`��4�Ē�ib�0��s�Ƒpa����&���j539.�f�,Ru� Env
�����2�3H�z�J9������h�Ф
Ҕ���2��2���� (K>L�n-TimФ������p�3�TS�����\kl�UTIL�"o���x�r "QMGl��!������1 "��S�T3�\kcmno��SФ�T2���ut�.�l�readc�}�exPY�ܤ�r��\��l�҄Фw�3��2C�*� -�C�D�E!Ĥ� .�4�C� R CV̴�҆��\p�Р���p�tbox��.�@��cycsL�:�RB�TE�veriOPTNE���;ӕӂk�e�ߦ�a�ߦ�h�g�ߥ�DPN��g�p.v��r�ptlit��0�4��te\cy���>�tmnu3`�r�����5UPDT�������駣���ite �� sw�to�,���oolB�F"�Y���Q��(q��gr3��䪒���"�䴁w������߳��s��������������lS���bx A"O�� ����l��`��P���A�l\t��� ��������	�Co�l�e!��R C ��r��&r �m;`��Chang�Lq�T1 �rcm3�"��
� 6���"����sPa7���"��22B2��2D4�57�� CC�FM�H��accda��Q�c' ��KÕ0���K!����m o!���,$Á��! "
����/�/����	�Y�,$��)�,$sk(����m rC%tS1,$�+��k1�%unc.�,$oñ�1��sub������1��cce �5/!&��-/?-W/i&vs�}/�%#�#�/��.C��/� C%
�@?  U �&+��F:qt�
pD�Ѓ D	 � U�:7�Dxmov.�P��DPvc\5Q�tfr@PeC_~UYgeobdtg_y[tu���P���PTUIt�P�Sx�_�^z�_��\var�_�\xy\�_�[pcl`c�P脆�P�Ue�Pgri�psuaoskuti����ovfinfpo}��o�j�b�P���Qud\�aX��Pc�\Rrp�Qnƅ�P�v�P)t�m#qƆ�P�v�a+ro�g�a��\Q�?a+rp#al?a{�{spa��@�P�u�Q�t�_TZp�0<�osipkag3r�o>vlclay(�:�t�pT�d�pu?a�c�A������KtKa�P䒏��qTf|rdm��{rin#r���As� �2���|s�PLd�v�tv��v�h�0��ystn* џ�y%t'�1�p��D�p�uϑ#�ul�@o�W6�92�siupdl�]�Fo�vr�on��`1L��z�`\�r���il3�$|l4��ǉ#q5 4FyB�Տg{�`���{�wcmס���wxf�er�UYtlk2�pp߿UYconv��sicnv�Qʯx�ag��H�Z�lct�`ao�=�p��׭nit0믁�3�������  �� ?v	�v	$��alϑpm�r&�B�eWa���f�%�� ����I��߬�u�ͬ�KamT�f���c��w��roǁ#�5�����?� sm��y�a��y� ��������`����͐ϑ��p��m�Wa� 1���A�6�S�e�X� �ψ�\Q}��������� ��ĥw߉�西߭�� �߮�#q0��rs�ew����1�a��z긱n�@�.�۲;�d�������  � �Ad	T$�1 �p! P��e �Ne 	lf@C��@�s/�  ?�����8�� �������r�eg.�C=��o�99 ~@�����$FEAT_�INDEX  �z ���e� ILECO�MP :��=�1!!z�$#SETUP2 �;1%;"��  N f!$#_A�P2BCK 1<~1)  �)��/�/  %�/�/e4 �/�/>%�/$?�/ H?�/U?~??�?1?�? �?g?�?�? O2O�?VO �?zO�OO�O?O�OcO �O
_�O._�OR_d_�O �__�_�_M_�_q_o o�_<o�_`o�_mo�o %o�oIo�o�oo�o 8J�on�o��3 �W�{�"��F� �j�|����/�ď֏ e������0���T�� x������=�ҟa��� ���,���P�b�񟆯 �����K��o���� �:�ɯ^�����#� ��G�ܿ�}�ϡ�6� H�׿l�����ϝ���t@)t Px/ 2� *.VR��߅�*�@߂�F�j�T���PCrߛ߅�F'R6:����V���z�T �!���K�� ��q�S�*.F�ߢ��	�Ӑ���x^����STM ��'���S����iPendant? PanelS���HI���9���U�������GIF0;�p�������JPG���;��]oR�
�ARGNAME.SDTy�>�\"����Rc	P�ANEL1Y�%�>��e�w��2 �A/�//���/�3_/�/��/p/�/?�4�/I?�7?�/?��?TPEINS�.XML�?>:\��?t?�1Custo�m Toolba�r�?Q�PASS�WORDg?w�F�RS:\:O�? %�Passwor�d Config {OR��OSO�O�O��_ �OB_T_�Ox__�_�_ =_�_a_�_�_�_,o�_ Po�_Io�oo�o9o�o �ooo�o(:�o^ �o�#�G�k ���6��Z�l�� �����ƏU��y�� ����D�ӏh���a��� -�Q��������� @�R��v����)�;� Я_������*���N� ݯr������7�̿޿ m�ϑ�&ϵ�ǿ\�� ���y϶�E���i��� ߟ�4���X�j��ώ� ߲�A�S���w��� �B���f��ߊ��+� ��O���������>� ����t����'����� ]�����(��L�� p��5�Yk  �$�Z�~ ��C�g�/ �2/�V/���// �/?/�/�/u/
?�/.? @?�/d?�/�?�?)?�? M?�?q?�?O�?<O�? 5OrOO�O%O�O�O[O �OO_&_�OJ_�On_ �O_�_3_�_W_�_�_ �_"o�_FoXo�_|oo��o�o�`�$FIL�E_DGBCK �1<���`��� ( ��)
SUMMA�RY.DG�obl�MD:�o*n`�Diag Sum�mary+8j
C?ONSLOG �qn�=qCon�sole log��7kpMEMCHECK��2���qMemory� Data3�;g�� {)�HAD�OW(�����C��Shadow C?hanges���c�-��)	FTAP�����=��q�mment TB�D;�;g0<�)�ETHERNET�0�`n�q~���=qE�thernet ��pfigurat�ion��B`%�DCSVRF/��'�@��C�%� ve�rify all�C��c1p� �DIFF8��0�ůD��%Z�diffǯ{��q�1�������J� X�q�|�=	�CHGD�&�8�ͿD�ܯ������2Ŀ����R� `�yτ�GD�.�@����D�����FY�3�ϳ���Z� hρߌ�GD$�6�H����D�����UPDATES.$��
�ckFRS:\�"�c�>qUpda�tes List�c�`{PSRBWLOD.CM��blN����e��pPS_ROBOWEL\�6o+� =�loa��o����&��� J���n�����9�� Jo���"��X �|#�G�k �d�0�T�� �/�C/U/�y// �/�/>/�/b/�/�/�/ -?�/Q?�/b?�??�? :?�?�?p?O�?)O;O �?_O�?�OO|O�OHO �OlO�O_�O7_�O[_ m_�O�_ _�_�_V_�_ z_o�_oEo�_io�_ zo�o.o�oRo�o�o�o �oAS�ow� *��`���+� �O��s������8� ͏ߏn����'��� � ]�쏁������F�۟ j������5�ğY�k� �������B����x������C�үg�v���$FILE_N�P�R]���Y�������M�DONLY 1<���U� 
 � �ۿ(���L��5��� Y��}Ϗ�ϳ�B��� ��x�ߜ�1�C���g� �ϋ�ߘ���P���t� 	���?���c�u�� ��(����^����� ��$�M���q� ����� 6���Z�����%�� I[���2�����VISBCK�����ų*.VD��*� FR:\�V� Vis�ion VD fileVd��� ����	/./�R/ �v/�//�/;/�/_/ q/?�/*?<?�/`?�/ �??�?�?I?�?m?O O�?8O�?\O�?�?�O !O�O�O�O�O{O_�O !_F_�Oj_�O�_�_/_��_S_�_w_�_o~�M�R_GRP 1=LeC4 w B�`	 ���lo~li`۬B���D��f�nӺMT� ��� ����e `i`a�o�khb�h�o�d�cic.N����L�K���?M� �H>5gE��|��i`@4��B���Az�?��Bf��9�f��l}A��A���A�8A�?�A�y��pj{i`F@ �qhq�y��~g�fF6��D�MqD�� �BT��@����l}?pD��6����l���5���5��|�l}B����B�C�B��jZBj�ZB}x�BX�~�e9�B�B�(��A�}jA��cB�dl叐�A������A�܏e�P���t�  �@���@h0�?�\	@�B� �����Ο��+�� O�:�_���p�����veBH` �<ā��A`0O����'�d
��Z��WZ�l�/�FX
��A@���@�33;@����\��[���ѿ�z��񿋯� *��N�9�r�]ϖρ��<�G�=��<�m]<�+�=~�m<c^���8eN7����7ѷ7�wx7;��51��Ϡ	ߤ��?߾d2^`Y�b`�b`�����TF�`Үb` b`�0�����C�^o�� �o�o�߸o��o��  ]�(߁�l������ ������#��G�2�k� V�{������������� ��1 ��- �)������ �0T?xc� ������/') �'/M/_/q/8��/�/ /�/�/�/�/?#?
? G?2?k?V?�?z?�?�? �?�?�?O�?1OOUO @ORO�OvO�O�O�O�O ��_��J����`_*� �_N�_�O�_�_�_�_ oo'oMo8oqo\o�o �o�o�o�o�o�o�o 7"[Fjh� x�t��!��E� 0�B�{�f�����Ï�� �ҏ����A�,�e� ,/���������/�J� ���=�$�a�H�Z� ��������߯ʯ�� �9�$�]�H���l��� ��ɿ��ƿ���#��O �OV� _z�D_V_��z_ �Ϟ_���
�C�.� g�Rߋ�vߛ��߬��� ��	���-��Q�<�N� ��r������� ��)��M�8�q�\��� �������������� 7"[Fk�|� |����֟3� WBg�t��� ��/�///S/>/ w/b/�/�/�/�/�/�/ �/??=?(?:?s?:� LϦ?p��?�Ϧ� O�� $O��T?]OHOZO�O~O �O�O�O�O�O�O_5_  _Y_D_}_h_�_�_�_ �_�_�_�_o��@o
� go*owo�o�o�o�o�o �o	�o-*cN �r������ �)�;�M����� ����ˏݏď��%� �I�4�F��j����� ǟ���֟��!��E� 0�i�T���x���ï�? �?��O��?OO� t�>O������ѿ��ο ��+��O�:�s�^� �ϩϔ��ϸ������  �9�$�6�o�6o��Zo ��R����������5�  �Y�D�}�h���� ���������
�C�U� �y�����d�����:� ����+Q8u `������� ;&_Jo� �����//گ 4/��x�j/4��/X�n/ |��/��/�/!??E? 0?B?{?f?�?�?�?�? �?�?�?OOAO,OeO PO�OtO�O�O���O�O _�O+__O_:___�_ p_�_�_�_�_�_�_o  ooKo6oooZo�oZ� �o�o�o�o��xo
 G2kR���� �����1��.� g�R���v�����ӏ�� �	��-��Q�/*/ ��N/��r/�/ޟ�/� �/)�D�M�8�q�\��� ���������گ��� 7�"�[�F�k���|��� ��ٿĿ���O�O�O�� W�B�{�fϟϊ��Ϯ� ��������A�,�e� P߉�t߆߿ߪ��ߪo ��+�=�a��߅� p�����������  �9�$�]�H���l��� ������������#�G2W}h�p���$FNO �����_�
F0� � } #�1 D|��� RM_CHKT_YP  � �q��� �� ��O=M� _MIN� m�����  �X� SSB_CF�G >� ~�Jl�A�j|�TP_DEF_OW  m����IRCOM�� ��$GENO�VRD_DO�����THR �d�d�_ENB�� �RAVC_GRP 1?3� X�e/��/ �/�/�/�/�/�/�/?  ?=?$?6?s?Z?�?~? �?�?�?�?�?O'OO KO2OoO�OhO�O�O�Op�O�O�O�ROU? �E� q�������8�?�#�O__K_m_o_ꐖ  D3���_Ed�_q�@A��\Bȡ���R��>Y_6 SMT
<#FC-�Ufoxo�o��HOSTC,1�GY?��_ 5	�h�k�o�f�oyeCU gy�z1�������p	anonymous�5�G� Y�k�w��o�o�o��� ���*�<��`� r�������ˏ	��� ��&�8��������� �����ȯگ���M� �4�F�X�j�����ݟ ��Ŀֿ���I�[�m� ρ�fϵ��ϜϮ��� ��}�����,�O�P� ��t߆ߘߪ߼��� /�A�C�(�w�L�^�p� ����ϸ�������� ��a�6�H�Z�l�~��� ��������9�  2DV��z��� ���#��
.@ ������������� ��//g</N/`/ r/�/����/�/�/ ?Qcu��/[?� �?�?�?�?�?)/�?O "O4OFOi?�/�/�O�O�O�O9m�aENT {1H[ P!^O._  `_?_ ._c_&_�_J_�_n_�_ �_�_o�_)o�_Moo qo4o�oXojo�o�o�o �o�o7�om0 �T�x���� �3��W��{�>��� b���Տ��������� A��e�(�:���^������㟦�QUIC�C0�̟ޟ?��1 @��.����2��l��~�߯!ROUT�ER௼�ί/�!�PCJOG0���!192.16?8.0.10	��GNAME !�J!ROBOT����NS_CFG 1�G�I ��Auto-st�arted/4FTP:?�Q?SOB� �?f�xϊϜϮ��?�� �����+�߿�P�b� t߆ߘ�6����� (�J� �1�C�U�g�6� ����������x�	� �-�?�Q�c� ?2?D? ���������) ��M_q����: ���%t��� ��m������� ���!/3/E/W/z {//�/�/�/�/�/6 HZ ?n/S?�w?�? �?�?�?�/�?�?OO <?=O�?aOsO�O�O�O �/
??.?0O_d?9_ K_]_o_�_PO�_�_�_ �_�O�_�_#o5oGoYo ko�O�O�O�O�_�o&_ �o1Cogy ����oT��	� �-�|o�o�o�o��� �o��Ϗ����)� ;�M�_�q���������˟ݟ�ÿT_ER�R I�����P�DUSIZ  j�^���$�>=�?WRD ?޵w���  guest+�}������ůׯ��SCD_�GROUP 2J�� �`�1���!��L_����  ��!�	 i�-	�E����Q�E EATSW�ILIBk�+��S�T 4��@��1��L�FR�S:аTTP_A�UTH 1K�<�!iPenda�n������!�KAREL:*8���	�KC�.��@��VISION SET���u���!�ϣ�������� 	��P�'�9߆�]�o����CTRL L���؃�
��FFF9E3���u���DEFAU�LT��FAN�UC Web S_erver��
�� e�w���j�|��������WR_CON�FIG MY��X����ID�L_CPU_PC����B�x�6��;BH�MIN'��~;�GNR_IO��K���"��NPT_�SIM_DOl��v�TPMODNT�OLl� ��_PR�TY��6��OLN/K 1N�ذ��� 2DVh��M/ASTEk�s�w�}OñO_CFG�Ƙ	UO����CY�CLE���_A�SG 1O��ձ
 j+=Oas �������/�/r�NUMJ�x �J�� IPCH��x��RTRY_C�N�n� ��SCR�N_UPDJ����b$� �� �P��A��/���$J2�3_DSP_EN�~��p�� OBP�ROC�#���	JO�G�1Q� @���d8�?�� +S? /?)3POS�RE?y�KANJI_� Kl��3��#�R�����5�?�5C�L_LF�;"^/�0EYLOGGIN� �q��K1$��$�LANGUAGE� X�6�� ,vA�LG�"S�߀�+����x��i��@�<𬄐'0u8������MC:\�RSCH\00\���S@N_DISP T�t�w�K�I���LOC��-�Dz�U�=#�J�8@BOOK U	L0��`d���d�d��PXY��_�_�_�_�_ nmh%i��	kU�Yr��UhozoLRG_BU�FF 1V��|o2s��o�R���oq� �o�o#,YPb �����������(�U��D/0DC�S Xu] =���"lao����ˏݏ��3n�IO 1Y�	 �/,���� ,�<�N�`�t������� ��̟ޟ���&�8� L�\�n���������ȯ�ܯ�Ee�TM  [d�(�:�L�^� p���������ʿܿ�  ��$�6�H�Z�l�~�p�Ϣύd�SEV� �]�TYP��$���)߄m�1RS�K�!O�c�"FL 1Z�� ����߯����������	�:�TP�5@���A]NG�NAM�$�E��k�UPS PGI|%�1�%}x�_LOAD0�G %Z%CAL_TC� ����MAXUALRM ;'�I(��~���#� QV�#a��CQ[x�@8��n��"�1060\	 �F�	�Ϣ��� ���������� D '9ze���� ����R= va������ ��*//N/9/r/�/ g/�/�/�/�/�/?�/ &??J?\???�?k?�? �?�?�?�?�?�?"O4O OXOCO|O_OqO�O�O �O�O�O_�O0__T_ 7_I_�_u_�_�_�_�_��_o�_,o��D_L?DXDISAc����MEMO_AP�]�E ?��
 �5i�o�o�o�o��o�o�o��ISCw 1]�� �o Td��\no�� �������I� 4�m��f���$����� ����!��E�ƏT� f�:�����ß����� z��ܟA�,�e�w�^� �����~������  �=���L�^�2����� ����߿�r� �Կ9��$�]�o�(t_MST�R ^�͂�SC/D 1_xm�W��� S�������=�(�:� s�^ߗ߂߻ߦ����� ��� �9�$�]�H�� l������������ #��G�2�W�}�h��� ������������
 C.gR�v�� ���	�-Q <u`r���� ��//'/M/8/q/�\/�/�/�/�/�/s�MKCFG `����/��LTARMu_2a��2� �#\`Y>G`M�ETPUT`�"�����NDSP_CMNTs506�5��' b���>�"1��?�4�5POSCFz�7�>PRPM�?��8PSTOL 1�c2}4@p<#�
aA�!aEqOG]OO �O�O�O�O�O_�O�O A_#_5_w_Y_k_�_�_�_�_�Q�1SING_CHK  +O�$MODAQ73d�
?�7:eDEV �	��	MC:>MlHSIZEs0����eTASK �%��%$1234?56789 �o�e�gTRIG 1en�� l��%��?   A$�Üf�YP�a,u��cE�M_INF 1f�>7 `�)AT&FV0�E0N�})�qE�0V1&A3&B�1&D2&S0&�C1S0=�})GATZ�� �H� E��q9m��xAu��� X�������� �� ����v�)���я ��П�������*�� N�����7�I�[�̯ ן���9�&���\� ���g�����i�ڿ�� ����ï4��XϏ�i� ��A���m�������� ��ѿB����ϊߜ� O������ߟߩ���� >�%�b�t�'ߘ�K�]� o߁�����(�_�L� ��p�+����������.�ONITOR�0G� ?ak   	?EXEC1�#U2345T�`789�#��xxx *x6xBxNx@Zxfxrx2U2�2�2�2�U2�2�2�2�U2�33�3�aR_GRP_SOV 1g�y�a(�Q�>�9�?�h����?��<���@�,Ѯ�Hm�a_Di�n�!P�L_NAME �!�5
 �!D�efault P�ersonali�ty (from� FD) �$RR�2� 1h)de�X)dh�
!�1X d�/d/v/�/�/�/ �/�/�/�/??*?<? N?`?r?�?�?�?�?�?�82S/�?O O2ODO@VOhOzO�O�Ob<�? �O�O�O�O_"_4_F_�X_j_|_�_LhR� �1m)9`\b0� �_pb�Q �@D�  �Q?���S�Q?`�QaAI?�Ez  a@o�g;�	l�R	 O0`4b@4c�.a�P�Jd�Jd�K�i�K�J����J��J�4�J~��j0Ea�o-a�@��o�l�[`@�z�b�f�@�S��a�Q�o��c�=�N��
������T;?f�
���m[`��*  �p  ��$p> p�$p���o?��?�����	��o�Bntr�Q�s�kse�}�l�p��  �pu`j7  #p��vks��� 	'� �� �I� �  ���}�:�È6�È=����N��b@�^�d��n�Q���{�RȒx���nN. ��  �'���a�`@a��@�t�@p@hp�n[`CpC0��f0�+pB/pC3}��P�@%�Ea�  oo�$|m����gA%���. ���z!�`�P���QDe����˟��(��m��� �t O�� ru �4 �R�c��sO� :�u�a�P~�` �?�ffd��!�����7� ���گ쬛af��>搠���iP�P;�e�0S�_�c���>LX��s��b<	�I<g��<#�
<2���<D��<��a
vo��¯�S��S|.���?fff?u��?&찗d@T����?�`?U��?X����Z� ��T:z�TB��Wa�з *dů�ρϺϥ����� ���&�8�#�\�h�+�F. Kߘ�G߼�3����Wɯ���G�@ G����X�C� |�g�y��������� �jZ���ￏQ��� �ߙ�����3����� ��/A��t_�(��������� �d���@+FpA�IP�t��%���[`B�0�����<ze�cb!@�I�
�M`B@���@`�9@y��?�h�� �@�3�[�N��N�N�E?��<�/:/L ��>��ڟ�A��p�C�F@�S�b/DpX������@�t�?�%�h��`/q�G��Gkn�F&�Fצp�E,8{�/ F��ZG���F��nE�DE�,ڏ�/� ����G��F7��F��ED��.� �C?.?g?R?d?�?�? �?�?�?�?	O�?O?O *OcONO�OrO�O�O�O �O�O_�O)__M_8_ q_\_�_�_�_�_�_�_ �_o�_7o"o4omoXo �o|o�o�o�o�o�o �o3WB{f� �������� A�,�Q�w�b������� ���Ώ���=�(�@a�L���p�����(r!�3�ji��r���<ꕢ�3Ա�ڟ�y�4 ����y���P�2�D�&��jb^�p�1w���������ʯ����ܯ� �s�P^�PD�c�`�m���y�\������Ӱ�¿Կ� ����.�G���� }ϳϡ���홍�U�_�J���$�y.�@�v� d�z߈ߚ�x�4����@���� ��D�.�2� ;�$[�G�[�^��B���B��CH � ^����u����������p�h�M�_��q����������"^�^�Y�m�2��
 ����#5 GYk}����p��h*�� ��>��x}��$MS�KCFMAP  ���� �����m�N"ON�REL  6��9_�"EXCFENBk
7]��FNC�}JOG_OVLIMkdu�yd"KEYk��"RUN���"SFSPD�TYU��v_SI�GNk}T1MO�T�z"_CE_GRP 1n��9\���/���/ �/4��/?�/2?�/'? h??�?C?�?�?y?�? �?�?O�?@ORO	OvO -OoO�OcO�O�O�O_��O*_<_#_`_-�"T�COM_CFG 1o/���_�_�_}
|Q_ARC_��6��UAP_C�PL�_�NOCH�ECK ?/ 5�;h9oKo]o oo�o�o�o�o�o�o�o��o#5GTNO_WAIT_LF'l5y"NT�Qp/z���q_ERR�!s2q/_�� R_���"�:�L�^dT_MO�sr�}, ��P_��_�_PARAM�rs/������MW���� =e�345678901.�@�R� )�q���_�����˟��0��ݛLW�3�E��؏i�cUM_RSPACE,��������$ODRDSP��SI&�OFFSE?T_CARToݨ�DIS�ݢPEN_FILE�I!�Q��v�POPTION�_IO���PWO_RK t�'�C T�|�C�������䖱Z���	 ��m���A����i�_D?SBL  ��v����ޡRIEN�TTOj��C����8=#�?�UT�_SIM_DJ��6	��VàLCT u�}�����Q��>W�_PEXE���RAT���� ��>�UP ve�����������*�8���$��2�#h)d�eX)dh�O�X dY�ߑߣ� �����������!�3� E�W�i�{������������2n��)�;� M�_�q�����������<�����+= Oas���X���� O��1m(��O�(�.�g��"0 �дu� � @D�  �?���?р��D4  EzZ3�;�	l	 '0ӀS@SM�� �i�i �H)�!H,�H�8�Hm�G�?	{G�8��6��MV��� �C�)���)�����Ճ�*  �p � � > � # ��/$"�,���B,�Btr�«{���¼�/���/�"�# �,�0 �� �  �� ߽pj   ��&X�?MU	'� � 12�I� �  ����-=���8U?g;/�@}?�0 ~.ѱ�?;Ѳ���&H[N �?A'M�D,�> C)�f)�" B& �"O4B+�:�Q��@D1�o�o$����JWAD0�J@�A: �1�E &?�O�O#__G_2]��� �t �O� ru �4 ��R<�U��� :�%Ё�р� �?�fAf��@[�_�_V_{��o~��18р"o0j>�P�Q6YPрZo�W�rAdS�%�>L�w0�#�<	�I<�g�<5�<2���<D��<��`��l�_�ѳ|Mb�@?fff?�0�?&p:T@T��q?�`?U��?X�-q�iyB q5Ya��g I�_������ !��E�W�B�{���d� ����ՏLnpΏ/�~ʈG�@ G�� U�ȏy�d�������ӟ �������yB=� � �?p���/򏸯�߯ R���'�9��oN�`������~�����ۿƿ�B�ĮD�e�ֿ;�xҿ_�J�?��h�PoϨϓϸ��D4��b!�_@���� ߧ�������%�@I��)�M`B@���@`�9@y���?�h	� ��@�3�[N���N�N�E��<��/Y�kЖ>���ڟ�A�p��C�F@�S����pX������@�t��%��h��߉!G���GknF&��FצpE,8�{�� F�Z�G���F�n�E�DE,ڏ���ૐ�G���F7��F��ED��Mf��b�M� ��q��������� ��(��8�^�I���m� ��������������$ H3lW�{� �����2 VAS�w��� ���/.//R/=/ v/a/�/�/�/�/�/�/ �/??<?'?`?K?p? �?�?�?�?�?�?O�? &OO#O\OGO�OkO�O�O�O�N(]�3�j�i�O�a��	U�E3�Ա��O_�a4 ��%_7_�a�Pq�Q_c_ERjb}_��_1w������]�Y�_�_o�_1o�l��P�bPcn~� ��o�O�o{_�o�oY�`��o�o,/; M#�f0o���� �Y�et�~�i#�1�C�yM�_��������� ��{bS�Ԏ��	�?�h-�c�Mj2���$�V'G�z}�B����B��CH�}�9� ֟�����0�B���wl�~�������Ư*�T���\�r�qQ��U
 ί �0�B�T�f�x����� ����ҿ���χ���� ��]{x}���$PARAM_MENU ?Յ��  �DEFPU�LSE�	WAITTMOUTl��RCV� �SHELL_WR�K.$CUR_S�TYLj���OsPT����PTB�����C��R_DECSNw�Te'�!�3�E� n�i�{ߍ߶߱������������F�A�US�E_PROG �%P�%B��V�CC�R��UeXÚ�_H�OST !P�!�����Tt`����Ŀ�����4���_T�IME�� �T�  �A�GDEBUG���P�V�GINP_�FLMSK]���T�R����PGA�� 2|�[���CH�����TYPEM�Y� A�;�Qzu��� ���
)R M_q����� ��/*/%/7/I/r/ m//�/�/�/�/�/?���WORD ?	>��	RS��C/PNS�E��>2sJO���BTE����TRACECT�L�PՅZ� }a` a`�{`�>q6DT QexՅ�0�0D��7���0��l�2�Sc�5{a�0��B ���7�0�2�0B�0B��0��2��2�4��4	�4�4�4��4�4�4 ��2��4�4�4�4��4�4�4�4(�4��2�4�4��*�2!�4"�4#�4��*�2&�4'��O&O 8OJO\OnO�O�O�O�O �O�O�O�O�4%X�1U(�4)�4*�4+�4U,�4-�4.�4/�40 _2_D_V_h_z_�_ �_�_�_�_�_�_
oo@.o@oRodovb�11�4U2�44�45�46�4U7�49�4:�4;�4U<�4=�4>�4?�4	@�4�9�o�o�o�o �o�o�o&8J \n������ ���"�4��1�= � 2�D�V�h�z������� ¯ԯ���
��.�@� R�d�v���������п �����*�<�N�`� rτϖϨϺ������� ��&�8�J�\�n߀� �ߤ߶���������� "�4�F�X�j�|��� ������������0� B�T�f�x��������� ������,>� bt������ �(:L^p ������� / /$/6/H/Z/l/~/�/ �/�/�/�/�/�/? ? 2?D?V?h?z?�?�?�? �?�?�?�?
OO.O@O ROdOvO�O�O�O�O�O �O�O__*_<_N_`_ r_�_�_�_�_�_�_�_ oo&o8oJo\ono�o V�o�o�o�o�o�o "4FXj|�� �������0� B�T�f�x��������� ҏ�����,�>�P� b�t���������Ο�� ���(�:�L�^�p� ��������ʯܯ� � �$�6�H�Z�l�~��� ����ƿؿ���� � 2�D�V�h�zόϞϰ�������$PGTR�ACELEN  ���  ��������_U�P y���2�������_CFG z�S������<��� <�Z�l�<�$��DEFSPD e{/��a������IN'�TRL �|/���8Lԃ�I�PE_CONFI�+�}��t�<�x�LID(��~/��GRP s1���������@�
=�[����A?C�C
��XC)��B�Y�r������dL��z������� 	� r�N��Ҩ�� #´����B�����������A���> �6>7�D_�������� ='�=)��������� 	B-��Q�Mx���  Dz����
��&L 7p[���� ��/�6/!/Z/���
V7.10b�eta1<�� �B=q�"`ff�@��">���ާ!=��͏!A>{ff�!@�ff�"��\)�"D��?�  �!@�!� �!Ap�#W��h/??*?<?K;�w����O/�?K/�?�?�?�? O�?O>O)ObOMO�O qO�O�O�O�O�O_�O (__L_7_p_[_m_�_ �_�_��_ o�_$oo !oZoEo~oio�o�o�o �o�o�o�o DQy<{/�#F@ {yw} �y{ջy�-��� ���/�Z?l?~?w��� t�����я������� ��O�:�s�^����� ����ߟ�ܟ� �9� $�]�H���l�~����_ ۯ�����5� �2� k�V���z�����׿¿ �����1�\n�j� |϶�������	� 4�F�X�j�c�χߙ� �߽ߨ��������)� �&�_�J��n��� ��������%��I� 4�m�X�����ί���� ������!E0B {f������ H�Zό�Vh�� �ϊ����� �2� D�V�O/�s/^/�/�/ �/�/�/�/�/? ?9? $?6?o?Z?�?~?�?�? �?�?�?O�?5O OYO DO}O�O���O�OtO�O �O_�O1__U_@_R_ �_v_�_�_�_�_�_" 4FxBo|��� �o��o�o//0/B/ ;�__J�n�� �����%��I� 4�F��j�����Ǐ�� �֏�!��E�0�i� �O^���N�ß՟���� ���A�,�e�P�b� ���������o o2o To.�hozo�o�����o ��Ϳ�o
گ'�֯ K�6�o�Zϓ�~Ϸ��� ���������5� �Y� D�Vߏ�z߳ߞ����� �����1��Uy� ��:���������	� ��-��Q�<�u�`�r� ���������� T�f�x�n����� �������7" [Fj���� ���!//E/0/i/ T/f/�/�/�/�/�/�/ ?�//?A?l�e?w?&? �?�?�?�?�?�?�?O O=O(OaOLO�OpO�O �O����*�O_@R�dZ_l_��$PL�ID_KNOW_�M  ����A�TSV ����P�[?�_�_o�O�&oo#o\o�B��SM_GRP 1��Z�� dI`�o�o$Cf�d����D��TPbj �oLk�f�o"~�U�o> n2T�~� ����7�4��� p�D���R���ʏ���� ������6�
�T��*�X�����QMR�c��m1T�EGQK? GR� �(�#���[��/�A� S������������$� ���W��+�=�O��� ��������� ����S�Ͻ�ST�a1 �1������P0� @����E�� ����������M�0� B�T�fߧߊߜ����� ������7��,�m���2�����A�<��z�3�������A4���������5)�;�M�_���6x���������7�����������8(:L��MA/D  ���� ���PARNUM � ��Ko���S+CH�
 �
�8�S+UPD���xaq{��_CMPa_�`� <Pz '�U~�ER_CHK�����Z���RqS���_�Q_MO� ��%_��_REWS_G����� � �v/{/�/�/�/�/�/ �/�/*??N?A?r?e?w?J'��W,g/�?L% ��?�?�?N#(��?O ON#w�4OSOXON#�� sO�O�ON# �O�O�O�N#d �O__N"V �1��Uua�@cX���Pp�P$@cW�،P��P@@cV���P�"THR_�INR���pbA%dޠVMASS�_ Z��WMN�_�SMON�_QUEUE Q��e��`Ȩ`�N�U�N�V�2`�END4a6/NiEX1E]oNeWBE\`>o>/cOPTIO;g?+�2`PROGRAM7 %j%1`O_��0bTASK_I���nOCFG �o�9pDATuAɓ�B{@ev2w������z� �+�=�O��s�����x����nzINFOɓ��}�!dr��!�3� E�W�i�{�������ß ՟�����/�A�S��e�w�҇ބ��| ��98q�DIT �Bׯj~WERF�L~hwS~�RGAD�J �ƪA� � ,�?E�8��Q�I�ORITY�W��>�MPDSP�a��j�U�WvT�OG��_TG���Rj���TOE�P1�ƫ� (!AF�PE�5 ���!tc�p��%�!ud|�?�!icm<��Q_��XY_<q��Ƭ�Oq)� *0������Op����� �������<�#�5�r� Yߖ�}ߺ��߳�������&�*�PORTT�a�OpA%��_CARTREP�~`ƭaQSKSTA��X!*SSAV`��ƪ	2500H809u�T毙䕣U�ƫ�����`�X#�$�6�m�URGeEU`B��A)WFP�#DO�V�2�W�q��?Q�WRUP_DELAY �Ư>e�R_HOT�hwR�%z����R_NORMAL�n��6SEMI:y�_QSKIP���X%;�x 	��� �����X%- ;%[mE�� �����!//E/ W/i///y/�/�/�/�/ �/�/?�/?A?S?e? +?�?w?�?�?�?�?�?�O�?+O=OOO1U�$�RBTIF��NaR�CVTM������m@DCR�����AB
�B}��>A��@��_ݧ������$�����V����HU���o���6��_ �<	�I<g��<#�
<2���<D��<��
+__{_�_)`���_ �_�_�_�_ oo$o6o HoZolo~oi_�o�o�o �o�o�o�o DV �_z������ �
��.�@�R�=v� a�����������׏ �*�mN�`�r����� ����̟ޟ����� 8�J�5�n�Y���}��� ȯ�����A�"�4�F� X�j�|�������Ŀֿ �ӯ���0�B�-�f� Qϊ�m��������� ��,�>�P�b�t߆� �ߪ߼ߧ�������� (�:�%�^�A����� �������� ��$�6� H�Z�l�~���{���� �������� 2V h������� �
.@R=O �s�����/ �*/</`/r/�/�/ �/�/�/�/�/??&?�28�AGN_ATC� 1��K �AT&FV0E�02;ATDP�/6/9/2/9�p8ATA2>,�AT%G1%�B960k9+�++�?,�1H�?,��AIO_TYPE'  EC/4?�REFPOS1 �1� K x�O[H/O/�O�M NO`O�O�O�O_�OC_��Og__d_�_+K2 1� KLON_�_o��_*o�_5A3 1� �_�_�_ o�o�o�o@oS4 1�Woio{o�o3W�oS5 1��o�oJ��|�jS6 1������]�H����S7 1��(�:�t���ݏ���S8 1�����Ϗ	���r����)�SMASK 1� O  
���ɗ'XNO�?���1.��8�1AMOTE  ��.DN�_CFG ��U���5�0BPL_RANGQ�K!Y��POWER ��Q5 a�SM_D�RYPRG %��%R���ȥTAR�T ����UME_PROׯ�d��.D_EXEC_E�NB  �5]�GSPD=����Y3��gTDB����RMÿ.��MT_ѐT��S��D0OBOT_N�AME ��S�;9OB_ORD_NUM ?���AH80�0I$�	��se	�\������ ��e��	@��}�D|��D0PC_TIMEOUT��{ xD0S232n��1�Q; L�TEACH PE�NDAN��j�5���=Q�x0Mai�ntenance ConsK"-���"+�t4KCL/)C�}�6��|�� No Us�e�=[߹�F���NPqO�ќ�5�_����CH_L@���U���	J��MAVAIL`���+���]�I�SPACE�1 2�=L �����p��扢�J@����8�? ��� ���V�w�N� �������������� 4�&G
l�}d	Q5 U1���������` 4&G
l}d�#��2������ ��2A/b/%/w/�//�/�3��� �	/�/-/O/^??B? �?�?�?�?�4�/�/ ??&?�?J?l?{O�O@_O�O�O�O�O�5�? OO1OCO�OgO�O�_��_|_�_�_�_o�6 _*_<_N_`_o�_�_ �o�o�o�o�o!�75oGoYoko}o+�o �o����)��>��8Rdv��H� ����ӏ%�F�-��[��G ��� R�;�
�� ����ԟ���
�� .�@����c���p���8�¯=�dؠ��ϟ�� �!�3�E�W�i�_�q� �����x��կ�� '�9�K�]�oρ�w��� ����Ͽѿ����5� G�Y�k�}ߏߡߗ���p������� `S� @��8堯F�"�*ل������ �������,���� V�h�2�<�N������� ������.L4 v�R\n�����
f�7�_MO�DE  ��MS ���&����AÏb��*	��&/�$CWORK_{AD]�5��!/R  ���t �+/^ _INTVA�L]���hR_O�PTION�& �h�$SCAN�_TIM\.�h��!R �(�3�0(�L8������!��3��1��/@>.?����S22�411d��8�1�1"3��@����?�?�?���IP���@���pJO\OnOE@D�� �O�O�O�O�O�O__�(_:_L_O���4X_�_�_��8�1��;�o�� 1���pc]�t���Di�1��  � lS2��15 17o Io[omoo�o�o�o�o �o�o�o!3EW i{����wc� ��	��-�?�Q�c� u���������Ϗ�� ��)�;�M�_��� `[����ğ֟���� �0�B�T�f�x����� ����ү�����$�7�  0��� om� �������ǿٿ��� �!�3�E�W�i�{ύ� �ϱ�������v��� /�A�S�e�w߉ߛ߭� ����������+�=� O�a�s�����ߖ� ���� ��$�6�H�Z� l�~������������� �� 2DVP�\�  �A����� ��%7I[ m�������/ �/C(/ N/`/r/�/�/�/�/�/�/�/?F;/?B?vF�x1 ;?�w=	12345�678{��l�@�P�?�?�?�?�?O9/2ODO VOhOzO�O�O�O�O�O �O-/
__._@_R_d_ v_�_�_�_�_�_�O�_ oo*o<oNo`oro�o �o�o�o�_�o�o &8J\n���o ������"�4� F�X�j�|������ď ֏�����0�B�T� f�����������ҟ� ����,�>�m�b�t� ��������ί����(��6yI�[�@��`���������Cz�  Bp*   ����254F��$�SCR_GRP �1�(�e@(�l��0�@ `1 �[1s	 )�3�C�<� t�vrY�8P�}�k�ܤ����95C����-u��ȡ����LR Mat�e 200iC Ə190�1Շ0LR2C �3�=OÆ��D�
f؜1u��2�U7��`1��v��@�u���	t�������h��$�^0�2� ��_2T�gϡϊ��o� F�D�f?��s���������ht ,Z�k`r�B�˰�P�N�g�rN�Aܰv�  @D���N�@����  ?� ��J�H˰��y�N�F@ F�`�� ����A,Qw b���n�N���`����B� �_J�n��� ��/�%//I/�΀E+:3��6?|?�5��
И/�/�#��@=�ò"�/pǢ� 3B�607�590@7����EL_DEFA�ULT  I��_�� ^1�MIPOWERFL  V�v5]2�0oWFDOk6 v5� �ERVENT �1���O�t3�C�L!DUM_�EIP?�8�j!AF_INEj0<O�$!FT�?=N�OaO!Q�O ��PO�O!RPC�_MAIN�O�H�8�O�O�CVIS�O�Iy��OE_!TP8P�PU<_�9d4_�_!�
PMON_PR'OXY�_�6e�_�_�XR�_�=f�_)o!RDM_SRV*or�9gouo!RR8d�o�4hdo�o!
�@�M�_�<i�o!?RLSYNC4y�8�oY!ROS�?�|�4H�tO �8c�����;� �_�&���J���n��� ���ȏڏ7�I���m�4���X����7ICE_KL ?%�;� (%SVCPRG1�����D!��3*�/��4R�DW��5z���6�����7ʯϯ�C��5�9��oG� ���o������D� ���l��񑔯�� ��7���_����� �4����]������ �����'��տO�� ��w��%ϟ��M��� �u���������� ?�A��Ͽ�ђ�؟� ����ɱ�������� ?�*�c�N��������� ��������); _J�n���� ��%I4m X�|����� /�3//W/i/T/�/ x/�/�/�/�/�/�/?�/??S?Ś_DEV� �9�M{C:[8�im4OUT_Rf1~6i8?REC 1���f0�0 f0 	� f0�2  
f0�4�1���3OMK�1�4=A%O^OAA���
 �Z�6 s;B�3AAqE@=�=A���2WG�1f0�)f0{f0U�Of2B>0�����/Q0A�O_�5��@��@�r�H�;@�  Ux�0}@U@��OK f0�f4�1af0��V_�2X0��@Ȋf0?�@�~_�__�U�2\�0��0��0��@����_ Rf0�f0�1=f0[f0��o�2T0��@̊f0*�@u*oco�_�eÆLH�0�0��R �  �RoTbmU�f0zf0�oT�2�Q��@�f06�@1z�ovo~K�L=A*�1(f0tf0�f0�_�c�f4e�=�ZZ Uf0k0��0Cf0�f0q��"~N@�LiI�1�2�f2Pf0Q>jI��zDf0f0�o.�g���φL"�f0i�0bf0��0�R�0V�b�f0f05/f0|~ 0��UE0��@�f0$�@PY�^�p���ՆL*�Ah�0=�Qpɀ��*b�ʈ�f0_^�f2�C0��@��A0����&��2\�AM��Up��A��p�Q<~��O��Ӧ�$2�,k�ҟ�2\&f0}��0�0Wf0�TZ��b�f0f0R~�)[���F��@ݒq0"ޯ�*�a@�� Z�H�~�l�������ؿ ������2� �V�D� zό�nϰϞ������� ����.��>�d�R߈� v߬ߚ���������� *��:�`�N��f�x� ����������&�8� �\�J�l�n������� ��������4"X Fh�p���� ��0B$fT��x�����5V� 1��<��`���A!O   -��P���a?_T�YPE�?k2HEL�L_CFG �4z:f2/ HL�/<7RSա�/�/�/ "??F?1?j?U?�?y? �?�?�?�?�?O�?0O�BOQK��p�!% QOO�O%��x�q�qQ��M�q�p�$�gBQ��d�O�O�&HK 1��+ �OE_@_ R_d_�_�_�_�_�_�_ �_�_oo*o<oeo`o�ro�oa&�#OMM ���/�o�"FTOV_ENM�t"!}*�OW_REG_U�I�o�"IMWAI�T�b���G${OUTrv$&yTIMuw��`VAL5>'s_UNIT�c�v�})MON_ALI�AS ?e�i ( he!� �� $�6�%��c�u����� D���Ϗ�����)� ;�M�_�q�������� ˟ݟ����%�7�� H�m������N�ǯٯ ������3�E�W�i� {�&�����ÿտ習� ��/�A��e�wω� �ϭ�X��������� ��=�O�a�s߅�0ߩ� �����ߊ����'�9� K���o�����b� �������#���G�Y� k�}���:��������� ��1CU y ����l��	 -�Qcu�2 ������/)/ ;/M/_/
/�/�/�/�/ �/v/�/??%?7?�/ [?m??�?<?�?�?�? �?�?�?!O3OEOWOiO O�O�O�O�O�O�O�O __/_�O@_e_w_�_ �_F_�_�_�_�_o�_ +o=oOoaosoo�o�o �o�o�o�o'9 �o]o���P�������s�$S�MON_DEFP�RO ����:� �*SYSTEM*  �l�*��RECALL ?�}:� ( �}�Bcopy md�:test_xy�.tp virt�:\output�\��over =�>1014497�28:951961  3�Џ⏻p�}7z���z.ls�~�������C�U��@z�z�����7�;�̟�ޟ�8��calpr��pc�2���D�V�����z���3��į֯�{��tcp@��%���H�Z�m�:���_dv�����5�ƿؿk�Fz������`��7�A�S�e�}9z�������4�����j�D ����ٜϵ�A�S�e� ������ϰ�3������i�tpdisc� 0=>lapt�op-3jv24�8ms:20980 �߬߾�O�a�t��tpconn 0 ��'�9������o�
xyzrate :������L��^�q�!���13960 �.�f������v����37224�448:8781�85 ��CU��A ���߄-<�d���5���_1��"�ASe�
2 #5�����ߑ� ��C/U/h�z�// 0/�/�/�/��
��/�" �/D?V?i{!0? �?�?�?�/
��?.?�?�QOcO�06�?��O  1O�O�OgO�?��&O �OI_[_n����_6_ �_�_lO�_�Π/�_DoVo�M?z��_"٠?<o �o�or��o&	�oEW�LE����"� ��w߉Ϩ,�D�V��C�ύݪo�� я��O?���/��O� a�t?�?��63�ğ֟ i�{������B�T�� ���/���ү�w����!���O�a���;�zRfrs:ord�erfil.da�t�dtmpback\/��6�ǿٿlz}2zTb:*.*��������P�b�pp��$SNPX_AS�G 1�������� P� 0 '%R[1]@1.?��?�ps%���Ͽ�  �����6��@�l�O� ��s߅��ߩ�������  ���V�9�`��o� ������������� @�#�5�v�Y������� ��������< `CU�y��� ���&	0\? �cu����� /�/F/)/P/|/_/ �/�/�/�/�/�/?�/ 0??%?f?I?p?�?? �?�?�?�?�? O,OO PO3OEO�OiO�O�O�O �O�O�O_�O _L_/_ p_S_e_�_�_�_�_�_  o�_�_6oo@oloOo �oso�o�o�o�o�o�o  V9`�o �������� @�#�5�v�Y������� Џ��ŏ���<�� `�C�U���y���̟�� �ӟ�&�	�0�\�?� ��c�u��������ϯ ���F�)�P�|�_��x�PARAM ���� ��	���P���p�OFT_KB_?CFG  �����״PIN_SIM  ��̶�/��A�ϰx�RVQST_P_DSB�̲�}Ϻ���SR ��	�� & CA�L_TCŵ�Ͻ��ԶTOP_ON_ERR  ������PTN �	��A���RING_PR�M�� ��VDT_GRP 1�����  	з��b� t߆ߘߪ߼������� �+�(�:�L�^�p�� ���������� �� $�6�H�Z�l�~����� ���������� 2 DV}z���� ���
C@R dv������ 	///*/</N/`/r/ �/�/�/�/�/�/�/? ?&?8?J?\?n?�?�? �?�?�?�?�?�?O"O 4O[OXOjO|O�O�O�O �O�O�O�O!__0_B_ T_f_x_�_�_�_�_�_ �_�_oo,o>oPobo to�o�o�o�o�o�o�o (:Lsp� ������ ���9�6�׳VPRG_�COUNT��8���d�ENB/�_��M��鴖�_UPD� 1�	�8  
M�������-�(� :�L�u�p��������� ʟܟ� ��$�M�H� Z�l���������ݯد ���%� �2�D�m�h� z�������¿Կ���� 
��E�@�R�dύψ� �Ϭ����������� *�<�e�`�r߄߭ߨ���������\�YSDOEBUGn�Ӏ� ��d��"�SP_PA�SSn�B?4�L�OG �΅ʹ� ���
�  ���� �
MC:�\`��a�_MPC f�΅����ҁ���� ҁ��SAV żi���� ����SV�TEM_TIME 1�΋W (J��F�{���%��T1SVGU�NSɀo�'������ASK_OPT�IONn�΅�������BCCFG �΋O� H�2!`;A�I�r]o ������� 8J5nY�}� ����/�4//�X/C/|/g/�/�/ � �,�/�/ ??�/�/H? 3?l?W?�?��?��0 �?�?�?O�?&OOJO 8OZO\OnO�O�O�O�O �O�O_�O _F_4_j_ X_�_|_�_�_�_�_�_ o�X�  o2oPoboto �_�o�o�o�o�o�o �o:(^L�p ����� ��$� �H�6�X�~�l����� Ə���؏�����D� 2�h�o������ԟ R�����.��R�d� v�D����������Я ����<�*�`�N��� r�������޿̿�� &��J�8�Z�\�nϤ� ����~������"�4� ��X�F�hߎ�|߲��� �ߤ�������B�0� R�T�f�������� ������>�,�b�P� ��t����������� ��(��@Rp�� �����$ 6ZH~l�� ����� //D/ 2/h/V/x/�/�/�/�/ �/�/
?�/??.?d? R?�?>�?�?�?�?�? r?OO(ONO<OrO�O �OdO�O�O�O�O_�O __&_\_J_�_n_�_ �_�_�_�_�_�_"oo Fo4ojoXozo|o�o�o �o�o�? 0BT �oxf����� ����>�,�b�P� r�t���������Ώ� �(��8�^�L���p� ����ʟ��ڟܟ�$� �H��o`�r������� 2�دƯ����2���P��$TBCSG_GRP 2����  ��P� 
 ?�  {���w�����տ ��ѿ���/�A�T�[���b�d0 ��p�?P�	 HBH�A�L�͌�@�B   C���϶ˀ���f��D����A���x���A��T$�9�ڧ6ff��f�@P�C��ώ�@�f߬��C��ߐ߮ߴޥ���%� �%�D�W�"�4����j�|�������?Y������	V3�.00s�	lr;2c��	*2�*�pO�A� ��ѳ33P�d��� x�J�y��  ������T�J�CFG ��el� o������������ =K
%�Kq\� ������� 7"[Fj�� �����!//E/ 0/i/T/f/�/�/�/�/ �/�/s���??(?�/ [?F?k?�?|?�?�?�? �?�?O!O3O�?WOBO {OfO�O�OP�<��O� �O�O�O0__T_B_x_ f_�_�_�_�_�_�_�_ oo>o,oNoPobo�o �o�o�o�o�o�o :(^L����� �h� ��$��H� 6�l�Z�|�����Ə�� ֏؏� ��D�V�h� z�4�������ҟԟ ��
�@�.�d�R��� v��������Я��� *��:�<�N���r��� ��̿���޿ �&�� >�P�b�ϒπϢϤ� ���������4�F�X� j�(ߎ�|߲ߠ����� ������B�0�f�T� ��x��������� ��,��P�>�t�b��� ������������ &(:p^��� �t�����6$ ZH~l���� ���/2/ /V/D/ z/�/�/�/j/�/�/�/ �/?.??R?@?v?d? �?�?�?�?�?�?�?O O<O*O`ONOpO�O�O �O�O�O�O_�O__ &_\_�t_�_�_B_�_ �_�_�_�_"ooFo4o jo|o�o�o^o�o�o�o �o�o0B�ox f������� ��>�,�b�P���t� ��������Ώ��(� �L�:�\���p����� ʟ��� ��_�*��_ �l�Z���~�����į �د� �2���h� V���z���¿Կ濠� 
�����.�d�Rψ� vϬϚ��Ͼ������ *��N�<�r�`߂߄� ���ߺ�������8� &�H�n�\���>��� ��x������4�"�X� F�|�j����������� ����
Tfx �D������ P>tb� ������// :/(/^/L/n/p/�/�/ �/�/�/ ?�/$?6?�� N?`?r??�?�?�?�? �?�?�? OODOVOhO zO8O�O�O�O�O�O�N�  PS �V$_R�$TBJ�OP_GRP 2���E�  ?�W<RCS��J\��@0�WP�R@T�P �� ��T�T ��Q[R	 �BL � �UCр D�*W[Q�_�_?fff~e:lB �P߆ff@`�33D  $a�U3o�>g�_�_po�l�P�e9�<�bbY��?�٪``$o�oUA�6�gD�`$�co�Q�uz9�P�A�a�P@a���C��Z`Ep�o]A6f�fpu`aD/�U�h�͔r��~�a�Rie Aq�`�q��@9q��|�d&`%���c3�33D�\P8����?�`?L�pAp[QB�b�k�}� ��z��� >�ffԁL����T�f��fo �� Nw@�*�8�f���r�,� ��П��ȟ��'�����F�`�J�X�����SC�Vء��	V�3.00�Slr2c�T*��TQ��� E����E�A E���E��3E�i�NE�!hE����Eۑ�E�I��E��E����E�rF��F�FM�(F�5F�BFaOF��\F"f,�z � E�@ E��� E�� E� � E����� E}����� EȆ��Ԏ�ᆰ� F�   F� F�$ Fj` F��@ F�P F��` 9�IR9��o���L�(_ ��V���LQ�8TESTPA�RS�XUP9SHR�k�ABLE 1ȒJ[4�SV�+� (�0�V�V�V�WTQV�	V�
V�V�T��QV�V�VȜ뱅�RDI��TQ��϶���������f�O n߀ۊߜ߮����ކ�	Sl�RS 0ړ��� ���������#�5�G� Y�k�}����������� ��/]k�o��*	�%� 7�I�����+�=�O����NUM  V�ETQ�PP� �밆�_CFGG ����Q@<P�IMEBF_TT�q��RS~�;VER��<Q;R 1=�J[
 8�R�P� �@5   ������// &/8/J/\/n/�/�/�/ �/�/�/#?�/?Y?4? F?\?j?|?{_�h�@R
<PMI_CWHANG R �3�DBGLVQ`I�R;Q�0ETHER_AD ?�E;@�S �?�?TO6V�0oROUTe!JZ�!�D�OwLSNM�ASK0HRSAA255.�E��O�O8T�OOLOFS_D�Iq��5IORQCTRL �s[���n]8]_�_�_�_ �_�_�_�_o"o4oFo��
�_Tofo�og�PE?_DETAIH3Z�PON_SVOF�F)_�cP_MON� �"P2�iS�TRTCHK ��J^mO�bVTCOMPAT�h;C�d��`FPROG �%JZ%  AL_�TCP=�n%QPL�AYr��j_INSWT_M�@ �|�g��tUSe]orLC�K��{QUICK�ME�0)�orSCR�EF�3Jtps��or�a�f��2�w�_{���ZyISR_GRP 1�JY_ ؛ 6 �����;�)�_�M��8����Y���� ���͕�����/�� S�A�w�e�������ѯ �������=�+�M��s�	12345G678����f�X`��1�Ћ
 �}�ipnl/۰gen.htm������0�B�X�Pa�nel setupF�}<�ϘϪϼ����� u�k��*� <�N�`�r��ϖ�ߺ� ��������ߝ�J� \�n�����I�?� �����"�4�F���j� �������������_� q�0BTfx�� ���� �>�bt�����3�~UALRM��pG ?J[
  �*/!/R/E/ v/i/�/�/�/�/�/�/��/??<?�SEV7  �n6�ECFG ��m��6��A�1   Bȩt
 =?�s3E �?�?�?OO+O=OOO@aOsO�O�Gz1ʂ��kC SΟ�OH7Isv?}{�`(%0?"_p _I_4_m_X_�_|_�_ �_�_�_�_o�_3o�L�� �M�OAoI_�E�HIST 1���i  ( �k`��%/SOF�TPART/GE�NLINK?cu�rrent=ed�itpage,,1 �q�`�o�o�'z�(�o�emenu�b955�`�ou���(:L148?,2 _XYd�`� ����}53�aZ������2�D���0n����"�4�À'LǏM~34�`�`4��������,K��nCAL�o��*�<�G�lY��`71�`MV��������í�)a�a)o ���%�7�I���ޯ s���������Ϳ\�� ��'�9�K�ڿoρ� �ϥϷ���X�j���� #�5�G�Y���}ߏߡ� ������f�����1� C�U����ߋ����� ����Я	��-�?�Q� c�u�x���������� ����);M_q  ������ �%7I[m �������!/ 3/E/W/i/{/�//�/ �/�/�/�/?��/?A? S?e?w?�?�?�/�?�? �?�?OO�?=OOOaO sO�O�O&O�O�O�O�O __'_�OK_]_o_�_ �_�_4_�_�_�_�_o #o�_GoYoko}o�o�o �oBo�o�o�o1 ?�ogy���� �o��	��-�?�� c�u���������L�^� ���)�;�M�܏q� ��������˟Z��� �%�7�I�؟���� ����ǯٯh����!��3�E�W�Bz�$UI�_PANEDAT�A 1�������  	��}/frh�/cgtp/wi�dedev.st�mc���ҿ����)�pri��.�Ip}�2�V�h�zόϞϰ� )���Ͻ������0� �T�;�xߊ�q߮ߕ���������Bv��� (� # Q�@�E�W�i�{� �������6������ �/�A���e�w�^��� ������������+ O6s�l�� ��������� 1C�g��� ����L	/// ?/&/c/u/\/�/�/�/ �/�/�/�/?�/;?M? ���?�?�?�?�?�? 0?Ot%O7OIO[OmO O�O�?�O�O�O�O�O _�O3__W_i_P_�_ t_�_�_�_�_Z?l?o /oAoSoeowo�_�o�o  O�o�o�o+�o O6s�l��� ����'�9� �]� D����_o�oɏۏ� ���#�v�G��ok�}� ������ş,����� ��C�U�<�y�`��� ����ӯ����ޯ�-� ����c�u��������� ��T���)�;�M� _�q�ؿ��|ϹϠ��� �������7�I�0�m� Tߑߣߊ���:�L��� �!�3�E�W��{��  ϱ����������r� /��S�e�L���p��� �������� =0$a����}�r� ����)�* ��Vhz��� �����.// R/9/v/�/o/�/�/�/��/�/?�������$�UI_PANEL�INK 1����  ��  ��}12�34567890 _?q?�?�?�?�?�4�� ]?�?�?OO1OCO�? gOyO�O�O�O�OYIY0�:�M��[0-/�SOFTPART�/GENA1?CO�NFIG=SIN�GLE&PRIM�=mainedit �OI_[_m_YJ_�$_M=wintpe,1@_�_�_�_XK  �_$o6oHoZolo oo�o�o�o�o�o�o �o
2DVhz �������� .�@�R�d�v��� ������Џ����M o0,M9P E=P�or?S�,Ico:�{�^�������˟ ݟ�����7��[�m�P������O���B0S0ߢ��C���/� %�7�I�[�m�`C��� ����Ϳ߿񿀿�'� 9�K�]�o��L���э� ��Q|���������� !ߨ�;�M�_�q߃ߕ� ��6���������%� ��I�[�m����2� ���������!�3��� W�i�{�������@��� ����/��Se w����.��� z�!E(W{ ^������/ �//A/���͡Ϸ�}� ���/�/�/�/�/?� 2?D?V?h?z?�??�? �?�?�?�?
OO�ϝ� ��dOvO�O�O�O�OE �O�O__*_<_N_�O r_�_�_�_�_�_[_�_ oo&o8oJo�_no�o �o�o�o�o�oio�o "4FX�o|�� ���e���0� B�T�f����/���� �����ُ���>�P� 3�t���i�����Ο�� O/�s/(��/L�^�p� ���������?ܯ� � �$�6�ůZ�l�~��� ����#O5OGO�� � 2�D�V�h���Ϟϰ� ������u�
��.�@� R�d�v�ߚ߬߾��� ���߃��*�<�N�`� r����������� ���&�8�J�\�n��� �������������m� "4ßXjM�q ������ BT7x����� �A��//,/>/P/ C�t/�/�/�/�/�/�/ o/??(?:?L?^?Ϳ ߿�?�?�?�?�? O O�?6OHOZOlO~O�O O�O�O�O�O�O_�O 2_D_V_h_z_�_�_-_ �_�_�_�_
oo�_@o Rodovo�o�o)o�o�o �o�o*�oN` r�����m ��&�8��\�n�Q� ��u���ȏ�������"���?�?�{��$�UI_POSTY�PE  �5_� 	k�{���_QUICKMEN  ��j������RESTORE� 1ו5?  ��/
�2�D�h�mc������� ¯ԯw���
��.�@� �d�v�������W��� ˿ݿO��*�<�N�`� τϖϨϺ����ρ� ��&�8�J���W�i� {��϶��������ߡ� "�4�F�X�j���� ������ߋ����y� +�T�f�x�����?��� ��������,>P bt����� �(�L^p ���I��� /�/��SCREܐ?��u1s]c-�u2M$3M$U4M$5M$6M$7M$y8M!��USER/ d4/F"T. O#ksW#��$4�$5�$6�$7�$8�!��NDO_�CFG ؜� � ,� ��PDA�TE �)�None V���SEUFRAME�  
��&,1R�TOL_ABRT87?��N3ENBX?I8?GRP 1�!��Cz  A��3 �1��?�?�?�?�?F!O"OG:ېUx81~g;MSK  {54�Ag;N41%a��B�%��O��VISCAND_MAXyE�I�c8�@FAI�L_IMGy@f����#�8�@IMRE/GNUMyG
�KRgSIZyC,���$�,SONTMOiUW0{D�%�VU��#�c�� �P�~�2FR:\�O� � MC{:\XS\LOG�V7B@4 !�O�_��Q�_o
�z �MCV�_�SU�D10fEX9k
��f�wV�2ۜ��p(ީ�=��͓o�� j�o�o�o�o�o�o�o  2DVhz���KPO64_?S��0��n6�uQ0L!I Q�z�x�qV� �|�f@�w�� =�	�xSZV�~�����wWAI��DS?TAT ܛ;�!@�_ď֏�$�����EP12DWP  ?��P G/����q�AP-��B_JMPERR 1ݜ��
  � 2345?678901��� ����ʟ��ϟ��$� �H�;�l�_�q����LT@MLOW���P�@μP_TI_X�('��@MPHASE � 53��CSoHIFTUB1~k
 <���Ob�� A�g���w���ֿ���� �����T�+�=ϊ� a�s��ϗϩ������ ��>��'�t�K�!��#�ޛ:	VSFT�1�sV�@M�� S�5��4 �0��U�A�  B8����Ќ�0p�����Ҫ��e@��ME*�{D�'q���q��&%�!��M�$�~k��9@��$~�TDINENDcXdHz�Ox@[O��aZ��S����yE����G����2�����������RELE�y?w�^_pVz�?_ACTIV���H<��0A ��K��B#&��RD�p��
1YBOX ��-�����2��D�190.0m.� 83��'254��2�p�&���robot�ԟ ?  pN g�pc� �{��v�x���$%ZWABC�3�=,{� 낆;-!/^/E/W/ i/{/�/�/�/�/�/?@�/6??/?l?!ZAT����