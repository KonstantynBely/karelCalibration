��   ��A��*SYST�EM*��V7.7�077 2/6�/2013 A�   ��	��BIN_CFG_�T   X 	�$ENTRIES�  $Q0FUP?NG1F1O�2F2OPz ?C�NETG  �D�NSS* 8 }7 ABLED? �$IFACE_�NUM? $DBG_LEVEL��OM_NAME �!� ETH_�FLTR.� �$�   ��FTP_CTR�L. @� LOsG_8	CMO>�$DNLD_F�ILTE� � SUBDIRCAP"n���HO��NT.� 4� H�ZA?DDRTYP� A =H� NGTHph���z +LSP� D $ROB�OTIG cPEEyR�� MASKa�MRU~OMGDsEVlFRDM*��DIS�BT�CPI�/ 3 $ARPSIZo�K_IPFpW_�MC-�F_IN�0FA~LASSܼ5HO_� IN{FO��TEL�G P�����R WORD  �$ACCE� L�V�$TIME�OUTuORT }�ICEUS� ���$O#  �����!��
��
�� VIRTUAL��/�!'0 �%�
���F����04+5�'�� =���!�!j?����; x?�5��=2~;#"SHA�R� 19 # Pf?O(4OHO 7OlO/O�OSO�OwO�O �O�O_�O2_�OV__ z_=_�_a_s_�_�_�_ �_o�_@ooovo9o �o]o�o�o�o�o�o <�o`#�G� k�����&�� J��n�1�C���g�ȏ ��쏯��ӏ�F�	� j�-���Q���u�����ן�ϟ0��7z _L�IST 1�=x/!1.k�09���j�1{��2551.��r����05i�2p���砖�����̯ަ3诂�_�� �2�D�ަ4`���װ��������ަ5ؿ��O����"�4�ަ6Pς���`vψϚϬ� �$��Q>�$% =��/5+5U�o!R��)���0H!� �����rj3_tpd���31 � �!!KC� �߿�(�'6��!C� ;���~��!CON� ������smond���