��   �A��*SYST�EM*��V7.7�077 2/6�/2013 A� ���$$CL�ASS  �S��(��D��D VIRTUAL%�7MNUFRAM�E AF�D� � 	� 88�?� ��}��y���� ��1=gQ s������	/��/?/��WNUM  ��>l�  �WTOOLa4� 
wN%M/  Bp�#C>3/U/�/1/�	?3????i?S>$�����D}?{:�1>�]�1ޣ1>Ӌ��&  G __?�?�?]?�? OO%OOO9O[O�OoO��O�Og,�!{&���&* 