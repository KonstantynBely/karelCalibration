��  /{�A��*SYST�EM*��V7.7�077 2/6�/2013 A�Q  �����ABSPOS_G�RP_T   � $PARAM  ����ALRM_RE�COV1   �$ALMOEN5B��]ONiI �M_IF1 D� $ENABL�E k LAST�_^  d�U��K}MAX� $LDEBUG@ � 
�GPCO�UPLED1 �$[PP_PRO?CES0 � ��1�FPCURE�Q1 � $�SOFT; T_I�D�TOTAL_�EQ� $,N�O/PS_SPI�_INDE��$�DX�SCREE�N_NAME {�SIGNj���&PK_F�I� 	$TH{KY�PANE7�  	$DUM�MY12� �3��4�GRG_S�TR1 � �$TIT�$I��1&�$�$T�$5&6&7&8&9'0''��%!'�%5'1?'1�I'1S'1]'2h"&��ASBN_C�FG1  8 �$CNV_JN�T_* �DATA�_CMNT�!$�FLAGSL*C�HECK��AT�_CELLSETUP  P� HOME_IO�� %:3MACR=OF2REPRO8�/DRUNCD�i2�SMp5H UTOB�ACKU0 �� �	DEVIC�#TIh�$D�FD�ST�0B� 3$INTERV�AL�DISP_�UNIT��0_D�O�6ERR�9FR�_Fa�ING�RES�!Y0Q_<�3t4C_WA�4�1�2HGX_D�#	� d $CARD_EXIST��$FSSB_T�YPi� CHKBoD_SE�5AGN �G� $SL?OT_NUMZ�AOPREV��G ��1_EDIT1
� � h1G=�H0S?@f%$EP<Y$OPc ��0LETE_O�KzBUS�P_CRyA$�4�FAZ0/LACIwY1KR��@k �1COMME=Ny@$DGV]Q@P� ���AL*�OU�B , !$�1V1AB0~ �OL�UR"2CAM9_;1 x�f?$ATTR��@�0ANN�@�IMG_HEIGHyA�cWIDTH�V�TCYU�0F_A�SPECyA$Mn@EXP;$� �Mf�CFcD X� $GR� � S�!1U`BfPNFLIxC`~d
UIREs3���AOMqWITSCH}cX`N.0S_d��SG0 � 
?$WARNM'@f���@� LI? �aN{ST� CORN�޴1FLTR�eTR�AT@0T�`  $ACC�1"p 8'|�'rORIkP�Cv�kRTq0_SF� ^4 �CHGI1 [ Tz`u3IPpTYVD�@*2 �P�`� 1zB*�HD�SJ* ��q2��v3�v4�v5�v6��v7�v8�v9�.:vqO�$ <� so��o�h�s1�PO_M�OR. t e0Ev�NG�8`TBA� 5c���A �����]@�����ϋP�0Ѕ*��h�`
P�@�2� �4,p�J,p_Rrrq�o@+�J/r/�J�JVq@�Cj��m�g��u6stP_}0OF� 2 w @� RO_�̿�WaIT8C��NOM_�0�1ەq3� ��cD �;���2�hP���mEXpG��0� F�p%r
$cTFx�JF�D3Ԑ�TO�3&@U=0�� ��H�24�T%1��E�� �e��f��f��0CPD�BG;a� k@$ƢPPU�3�f1):��A�AX 1�d�UN�$AI�3BU�FuF����! |��`��`PI�*�Pr�Mq�M~�����Fr�SIMQS@��G��QE�����[MC{� �$}1�JB�`S�}1DEC�������۵z� ���0CHNS_EMP�r$Gg�=Ǎ@�_��q3
p1_FP󔞡TCh�@`�b��@q0�c}�y�G�� V�A0Ԃ�!!���JR!0Ԃ?SEGFRA.pv �7aR�T_LIN�C��PVF������Y���Q���)B����( ' ���f�e�S���Q��.0��p�B��A����SI!ZC�ћ�z�T��g�������QRSINF 3��p����?�������؉���Lot��G�*�gCRC�eFCCC�` +���T�h��mh�SbA@��h�*�f��:�D�dd�c��C��PTA��`��w@�撀��EV���jF��_��F��N�&�G�� X�������1i��! ��,��hRGNP��0qF���R}�D���2}�LEWN��Hc6����C�K�vqRcDx :�L��ou2��ԊA6N`Co�$L	Gp��B�1aP��s@��dWaA?@���~0R���dME%`��d��_RAs3dAZ�C���z�OkqFC�RH`X`F�`��}��,�ADI;�  6b� ���`�p�`5c�n�S�@1�7a�AMP����PY8CU�M��CU��iQU� $�P��C�CG1�������DBPXW�O����p$SqK��2��DBT �TRL�1 ��Q0T�i� �P�DJ�4L?AY_CAL�1R !'PL	3&@�0�ED�Q5'�Q5'̡�!���1!�W�PR� 
�1 0Δ1" �PA$��q$�� �LB�)#�/�#mp�0$�/��$C�!%�/�$ENEqr�&�/�#d �REp�"'H ��O)@"$LF3#$�#xB� W;����FO[ _D0m�RO(@���u��j���3�RIGGER�6P�A%S���ETUR�N�2RcMR_��T�U�`?�u0EWM����GN�P��zB�LA��E��$$EP#�CP� ��&@D�Qk�C5D�mpD�A�#�p4\1i�FGO_oAWAY�2MO��tfQg�CS_7(<�QIS � ���c�C���A����B�t�Cn��A"�F9W���DNTV@��BVkQ�����S˳W�s�U�J&�U�� ��SAsFE�ZV_SV6b�EXCLUl���N��ONLA��SY���Q�tOTBa��HI�_V/M�PPLY�_�a��VRFY_�#�q�Bd�_ �)0���_+�Ip� �TSG3� *�b݀�0 AM��� a*����0��Vi.b>%fANNUN� r�LdIDp�U�2~S @�`mijarj�f�R�pOGI�"+��c$FOb�׀OT@�w1 $DUM�MY���d[!�d١��& �E, ` 8�HExs��b�S|B$�SUFFI��@ ��@�a5��g6�a��DMSW�E- 8��KEYI����TMZ1^ӌq�1�vIN����ir�. D��HOST? !�r���t[ `�t٠�tYp�pEM>����$��SBL��UL��/ �|3�����T50�!0 �� $9��ESAMP�ԕF���������I�0��$SUBe�Q�� �C�:��G�SAV��r���G�`C� ˇ�PnfP$80yE��YN_B�71 0��DIad�@�O���}$]�R�_I�� �ENOC2_ST � 2
�� J���L�q~S�`;����!3�M�I��1�:�p�4   L�3�M��0�0K�4<'a��AVER�q���}�M�DSP�v��PC�U���\ì�oVALUŗHE� ���M�IP@���OkPP7  �THS ����6�S�F�F�􁳠dL�0�T��SiC�Q�d:�ETo��5zrFULL_DUY�da�0��O�w��h�OT���0N_OAUTO�!6�pC$�\���cl�*
�C_��C����_��L�� 7/H *�L���n�b���$�0P�˴�� ֲ��[!���a��Yq��Tdq��7��8��9���0����1��1��1���1Ⱥ1պ1�1*�1��2
�2����U2��2��2Ⱥ2պU2�2�2��3
ʥ3��3����3��3�Ⱥ3պ3�3�3b��4
�����SE�"8 <��~��`�;�I�����/��QFE8�0�0� 9 ,��Q�? z@^ ?(�А��ER@#���Q�A��� :�`$�TP�$VARqI�<��UP2�P3; �pq�TD��S�|�1`3��� e�B;AC�< T�pr���)��bP�P o�IFI)�P ���U���P�& ��0��� =t ;'�Ԡ��P'�ST(&�� HR�&�r0E����	%�C��	���_Cr�N�r���B��p�h�FORC�EUP%bn�FLUS�`HN �E�h�^�RD_CMK@E(����IN_��&vP.g�REMM�F~Q��@M �� 3
K	9N0�EFF���N@IN�A��OVM�l	OVAl	TRO�V���DT��mDTMX���m{@�
���? �*[ ��CL��_:p']@$�-	_
�;_T��X
���@AQD� ���}��}!V1� R�Q��LIMIT_Ƚa椀�M��CLmd}�RIV	�a���EAR��IO*P�CC�����B�Bg�C�M@��R �GgCLF�G!DYM(�/�aR#5TWDGЍ�| s% �SS& �s> P�a�!r1���wP_�!�(�!1R��E�3�!3�+5�&O�GRA���?w�i�kPW��ONT��EBUG)S&2*��P{@a�_E @�:��Q�@�TER�MB5AK5��'ORIG0BK5���SM_�Pr�G0C\K5�P�TA�9D�6� �UPB�Eg� -zAa�@.P|Y3.@A$SEG�:vf ELEUUSE�@NFI,��2�1xޠp4�4B$UF6P�$�FQ4@�wAG0TQ�&�HSwNST PATm�<piBPTHJ�AߠE�p��2�P؀	E)��؁��1R�@�InaS�HFT_��1oA�H_�SHOR ܣ�6 ��0$�7�@Dq�'�O#VR#�na�@I�@��U�b �QAYLO=�z��I'"�oAj�!�j�ERV��:Qh� �J��OG @�B0����U�>���R!P"�AScYM.�"��1WJG�уES�A�YvR�U�T @���E)�ᥳEaP!�WP!�WOR @�MB��GRSMT�F�GR��3la�PA.@��`�q�uG� � ����T�OC�1�`P�@ �$OP��ဝpՓá� ��O��RE�`RC�AO�pтpBe�`RmE u�h�A���e$PWR�IM�ekRR_�c4��q.B H2H���p�_ADDR��H_LENGqByqnq�q��R��S�I H��S���q0Ӧu>Ӵu���u��SE�'�LryS��J $�<�`��_OFF��r�PRM� ��aTTP_�H��K (^pOBJ�?"ip��$��LE�`C!�ȠL � ��׬�AB_~T�S�s�S{`��*�LV�N�KR��eHIT���BG��LO�q t�fN�͂���`���`3SS{ ��HW��A��M�p`INC�PU�"VISIO �����+��t,��t,�~�� �IOLN���N̠�C��$�SLQb��PUTM_�$�`{�P x�V���F_AS�"O��$L��I���D�A��U�0�@Af��`q�<PHY���Ó�[���UO��#P `������ڔ� �2�pP���`(�L�p�Y�B� ��UJ��Q�z�NEWJO9G-G��DISx�[�1K-�f�#R 
�WA9V�ǢCTR�CǢ�FLAG�"[�LG�dS ���Y�3?LG_SIZo���`������FD)�I�4�E�*��D0� ��c$���𖶦����K���D0��� SCH�_��߅p�2�L�N��F�T���E �"~�������U
�
�r{`L�	�DAU/ŃEA�-��dE�;�G�H�bU�OGBO}O��Uh Aɒ���IT��y�[0ŖR;EC��SCR�𙃖ʑDIēS.@��RGO���˒����d��$����SU���W�Ĳ��Ľ�JGM$�MN�CH,�FNKEuY%�KM�PRGK��UFY�PY�FWDvY�HL��STPY��VY�@Y؀�Y�RS"��H1`uۺ�CT�� �R��� �$�U	�m�@��
R�ݠғ`�G=ن�@POd�ڻŦ�M��FOCUd�RG�EX��TUIK�I{�����	������I�M��@A�S�`��p�@������ANA����2�VAILl�C�L!�UDCS_H!I+4`�s_�Oe�
!"h�S���|�S����IGN4��F�J��9T�be�_BUj � �V !PT�$ *��rv�Ϥ&���a
�!W !Pi�'��T�0�1?2?3?�!��`� X � �i�=a�5���Ņ�IID� tbP5R�bOh X��\A�ST	�RF��Y� �@�  W$E�C�y�����_�� Y L �؟0��@���`q�Ftǀ�FwҬ�_ Z �p����b���>0C��[ ��p CLDP	��UTRQLI{��T����FLG�� 1�bO�D�����LD���ORG����� �hW>(�siT�r� 4\ �#0��վ�%Sy`T�70#0' ��$�!�#RCLMC��$B/T/�)Q��!=1I��p_d] d�R}Q73$DSTB�p`� �0!5��-8AX�R� /8I<EXCE�S�b 5Mp�1^��p2�Tt6��0_�p"6_A:&��;�G?Y80K�d` \��GROU��t$�MB �LI9�CREQUIRDB�aL=O#KDEBUr�1LYM��agbʑ`@h�C�"�1ND���`c`b���̨�CDC���IN'��C��Z`���H��N��a#�� t2�APST�� �c\rLOC�R!ITp��P�Ap��1�1ODAQ��d� X�ON�cF �R�fV�	X��b�U����u�FX0IG}G�� e �y @X�a��X�XR�Q%��Y	��X	��V<�0ғDATA$`�E�a��a�N��f t $MDEaI:�)Sf��^d�![g�H5P�@]ez��_cANSW�a^d�a��^eD�)BQz�� Xp�g �0CU4�V��`�=URR2{�h� D2�`A��A�! d$CALI&0ү�GS�w2K�RI�Nb�t<�NTEg�(i�bCu��=RBqg�_N�qjPukr����$ht�2kuyDIVF�&DHi0jp+�l �$Vp�C�$M�$Z0R<!T 0R����b�emH ?�$BELT˪Z_ACCEL���;�"�IRCO�݁m���T���$PSi0�L  ��U���Cp8��T�9�PAT!H���.���3]��Pl1_<�r��Ł�"S �Cr��_MG���$DD�9���$FW�`7`���.����DE�PPAB�Ne�ROTSPE!EՂ@L� JN�@�(0�]�$US�E_p�P&�ܦS�Y>��p�! �QYNr0A����OFFuan��MOU߁NGJ��܀OL~�ٔINC �d2Q��-2��� -2ENCSpa2U�X�+4R�IN�I]�0B����"n�VE��s>^�23_UPօp�/LOWL��[�` '���D>�2@Ep�]'��2C[pW�MOS���4MO��0�'PERCH  ��OV����蓼��� ���$�8S+�� 2@�������V�0^�O�L`�P��7O�U�UP"�8������TRK��AYLOA�J��1���]�͵³3P� �RcTI�1	�� MO� _�-2�28 �`4�w�ٳ��?�pDUM�2��S_BCKLSH_C]�P�ϐΦ ����bn�"�y�Ñ��!CLAL V��!8��� ��CHK �SՐRTY����C��
*!6a_�ä_U�M����C���SC�L�W�LMT_J'1_L< 0-օa:�E4�U�G�D�J�P�J�SPCd�ȑZ���&3�PC �3�H_A@d���C� cXT��.�CN_rN���".�S��%�V���@:����]�9���C' �SH�r�*�*! 9�9� p��^���9���3PA���_P��_�"�Ŷ�!ճ�����JG����~�OG|��,�TORQU��ON��޹*�B٢-�L*�L�_Wž�_�s�j��sj��sj�Ir�IJ��I�sFKP]�J�!X��c!�VC�0'42��1��{0��82���JRK��+� D�BL_SM���"Mζ@_DL�q�"GR�Vq�j�sj�sKH�_��I���
COS��LN- ��� ��p�	�p�	���ĺ�FZ� ٦KMY��D�TH�eT�HET0��NK2a3�s��s� CB�CB�sC&1n2���0��s��SB�s�N�GTS�1W�C.� 2Q�����$�'3$DU���8A!r �2P&�1Qb8V'$NE�4�PI� ��H�"%�v$�p�A��%�'���LPH�5�"h��"S��3� 33�"+3:2�pEV�(V�(�p�,V�*UV;V;V";V0;V>;VL9H�(�&�2P�-n�H;H;H";UH0;H>;HL9O�,�O�(O}I�.O�*O�;O;O";O0;O
>;O2F�"�Y��T�'SPBALA�NCE_T@SLE6�H_�SPHq��hR�hR3PFUL�ClX�R{W�R3Uz1=i
�UTO_�����T1T2�Y�2N ���`��Tq���Ps (d���T�O�p!�>L�INSEG����REVf��Q�DI�F��zy1j_g�r1k��OBUa��t$y�MI`���SLCHgWAR>��AB��~u$MECH��Tˑ�a��AX˱P�y��f�'�r�Pl 
p�bI��:�ROB��CR]�-u��#&��MSK_KP�tn� P �P_��R ��r_tn���18�c��a�_p`�y�_p�aIN�:a�MTCOM�_C���po  �݀g`4�$NO�RES��r��`�r7p 8U�GRJ��e�SD� ABג$?XYZ_DA�!F�r�DEBU:a�q����pq _P$��COD�� 1����`���$BUFIwNDXa�  !��MORRsr $�qU&���u��ӑy��^��bGi�s �� $SIMUL���8��>���F�OB�JEjP��ADJUySψAY_I���8�D���s�Ԑ_F-Iב=s�TZ�� c����`b�"�(�b`tp0G�D��FRIWÚd�Tg�RO%�A�Exb񊰓�OPWO> �Vpt0>�SYS�BU0[�$SOP���I�����U��b`PgRUN�rڕPArp�Dٖ�b��1�_OUbTΑ�a�t$�/IMAG��\pv �PDaIM��1�IN�[ �0�RGOVR!DY�˒���P�/�a�� L_�PB�}��¦�RB�� ��MLkᜪEDb��` �%N�@M��~���]��SLjPVpu x �$OVSLfS;DI��DEX���q �����o��Vb��N�A��'��,�'��D�M~Ҥ_SsETK�Vpv @U�^��ep�RI��j�
q�_�}�����Z�da|̀*� w H\q��`��ATUS<�$TRCx T�X�ѳ�BTMڷıI���P�4}Ѱ���Vpx �D\pE���β�0E�hbϱ�����ϱEXEհ����)�=��f�1ym�]p԰UP�L�s$�`6�XNN����������� �PGn�uzWUBñ��e��ñ��JMPW�AI[�P���LO�7��pFA`��$R�CVFAIL_Cwq�p��R9��p�c���(�}�"�-�AR_P=L��DBTB��,���pBWD ��pUM*�"�IG�7��Qc�GTNLW�"�}�Ry�iӻ�E�����^����DEFSP` G{ L\p�`��_��Ճ��UNI�����b��RD��Rb _LA`APͱ]����pUq|-��#��q�O��XPc�NN�PKET�
��Pq�Uq} h�ARSIZE����=���u�S̀OR��F�ORMAT�Pg�C�Oנq�<bEM�dL����UX��,�:���LIb�Uq~  �$�pP_SWI��`�� �/ G�b�A�L_ o���AR�rB���C�rD���$EL���C�_lі� � �c ���r��J30 ��r��TIA4Z�5:Z�6�rMOM��f��s���pB��A�Df��s����PU�NR����s������VF��Rt�� A$PI�&E�kqE� p-~-�-�W@C�0$��&�9q��gE��eSPEEDL@G�����Ծ�� ��)�9����)��	)���SAMWPx�08�1��MOVD�H$�_S`Y%nk%_��1�t�2�t����c�vd��8�H�PxIN� ��������(x�+(+GAMM<V|u!�$GETE��U�ٓD5�
�PL�IBRv���I�$HIu�_L�ݰpB�&�E�(A�.� �&LW�-�&�,�)	6�&1���f�`j��� $PDCK���ٓ_�����E��ီb7��a4��a9�� _$I��R�`�D�c�b~�Ե`LE@�qkq���81��0�Gq���`Vp�P/aUR_SCR��A�r���S_SAVE_�D��8Ex�NO5�C ��y�6�8@{$E�.{I ��G	{I�@�J�KP�q ��H� ���x"Ma o���s����d�@�6W2U�Cqy���M� �k�F�� aE��3�W<�@[�jQ!Wg@���U�R�R��ȥSc2jQM"��[CL��W��M)ATr� �� $PY����3$W`�fNG�O� `�b�b�b#�HЈ��a� ���c��X�O���Z�e��ހ�Rt� p䠰p�3 +zO�O�O�O�O�a5�_�r� |�E�8@ ��>vs�>v��8@_�kwVvy�Eހu%�!sB��\�P�"tP����PM&�QU5 �� 8*�QCOUܒ1 �QTH#pHO�L,�QHYS��ESe�qUE�p.BZ�]O��  q�P��̕%��UNְ�Q ���OE��p� P�2�3��AÔ�ROQG�����Q2(�O}��2������INFO�q� #�e����R�Ⱦ�OI��� (�0SLEQ�с��рi�C�{�D��L��D`� OK0r��!�E� NU!��AUyTTA�COPYqPu�?��`@ML�NI��M�X�Cᐛ� Y�R�GADJ�q�i�X�Q��$ഖ�`��W��P���0��������EX8�YC0b$�ѪObp�q���$�7_NA9!��������`��� �s Q���PORӸA�B�SRV0�)la�Y�DI��T_�� {�������������U5��6��7��8y�Ҿ�S8BL��m�MCS_F�p��PL9A8An�ȰR��9��Ѽ���$iB����d� �,�0FL-`L�C@Y�N�[�M��C?��GPWRc��L��!�ODELA��8Y5��AD�a��QSwKIP� �Q�Z4�OR`NT�Q ��P_4��ַ@lb Yp������ ����Ƞ��ՠ���������9�1�J2Rܻ L�� 4*�EXs TQ%����(Q�����p�����p���RD�Cf� �`��X9�R�p�����r��~A$RGEAR_� sIOT�2FLG��vi��M%PC��B�U�M_����J2TH�2N'�� 1������G8 T00 I�����MlѺ`I�\8AREFr1�q� l�h��ENA9B{�(cTPE�0� 1���i�m���^QB#���:��"������2�ҙ����������
&�3�Қ7�I�[�m�(��&�4�қ�����������&�5�Ҝ�1�C�U�g�y���&�6�ҝ����������
&�7�Ҟ+=Oa(s�&�8�ҟ������&�SMS�K�q�|��a��E�?A	��EMOT-EF����a@���(Q�IOQ5�Itc(P�POW�0L�� �pZ�����#p%�L��U�"$DSB_SIGN�1H)Q%���Cl�(P��/S232��b�i�DEVICEUS��,R'RPARIT|��D!OPBIT`Q�Y�OWCONT�R;�(Q��O'RCU�� MDSUXTAS�KT3N�p[0�$TA;TU`PV"�0RL����p_,PC9��$FREEFR�OMSp��%�GE�T�0�UPD(�A��2V"P� J���� !)$US�A^���6���ERcIO�P@bpRY�5:"_>@ �P}1�!�6'WRKI[D���6���aFRIEND<mQ�P$UFw����0TOOLFMY��t$LENGT�H_VTl�FIR��`-C�RSEN ;IU�FINR]��R�GI�1ӐAITI���4GXӱCI�FG2�7G1��Ѐ3�B�GcPR� A�O_~ +0!�1REЀ�E3�e�TC���Q�AVG �G8��"J���u1~! ��J�8�%���%m��5�0G4��X _0)�L|�T�3H6��8���%r4E3%GU�W�P�W�R�TD����T��а��Q��Tm�$V 2!����1���91�8�0U2�;2/k3�;3�: iva�9=i�aa�^SL�jR$V��SBV�E�V'�V�BK���� �&c�p��F�"{�@��2q�PS�E0��$.rRC��o$AŠFwPR��Gv]U�c1S'�� 7�QA6I�G� 0�@qV`��p�d`���E0�@��=��
B5S!� �"�aRg����R�6�MN AX�!$�A�0�L(A���rTHIC´1Y���h�t1TF�EI��q�uIF_C	H�3�qI�G�a�pG1bxf���m���S@���_JF��PR��ֱ�S��Ԁ�Od �$SР�Z��GROU�̃TO�T�t̃DSP�JcOG���#��_P㱂�"O�����j��&KEP(�IR����@�M�R@�AP�Qn�Ep^�`�!�[�SYS6��"[�PGu�BRKP�B �.��pIq�p`��M���΂�`AD�!<̃9�BSOC׆��NӕDUMMY1�4�p@SV�PDE�_OP�#SFSP_D_OVR=���1C���OR�C�Nm0�F.����OV��SFR��pU���Fn��!#��C��A�"�LCH����РOV(�s0��W�@M��ĥF:�RO�#ߑ�_�p��� @@�u@VE�R�ps0OFSu@CV? �2WD6���2��ߑj2Y���TR�!|���E_FDOY��MB_CM�D�B�BL�b>�f��att�V"Q�240/p��N�Gg�z�AMx�Z�0���¿_M~��"7�����8$CA�7�D:����HBK81��IO�5���QPPA�=�"�M�5��͵���DVC_DBxC~� �3"�Т�!"��1��糖�3��� �pН�*��U�3��CAB��2VӆP�ѣIP��c�O��UX~�SUBCPU�r	�S�P P���90^S�Q׹c��."��$HW_C�Т��S��c�A�A�pl$UNI�T��l��ATTR�I"���	�CYCL���NECA��J�F�LTR_2_FI`_�G(��9&�1LP��?�>�_SCT�CF�_��F_��6��FqS8!����CHA�1��wᇲ�"v�RSD��4"����q�_T���PRO��>�� E%My_ܠ��8d��a� d��a��DI�b0!�RAILAC4��9RM��LOÐ C��Q*q��3q���+PR��SQ�pU��Cr�s 	�FUN9C��@rRIN'P�0�0��u��!RA��B� ����F�Ğ�W3AR~���BLQ�����A��������DA`����	����LD)0 ��Q1�q��*q1�TI2rQǁ�p$�xPRIA1�"AF
B�P�!|ߠ�<`8�R���MOI��A��DF_&@��51��L�M��FA�@HRD]Y�4ORG6 H����A�0 �MULS�E&@"�Q��a ��G�	�����$�d$�1$1� ���0���� xm�EG�̃�`cARހ��09�2�o��z�AXE�RKOB�W�A��_��œSY������SN�WRI�@s1���STR�� ��(�E�� 	%1��AB( �/&�a�ӰkOT0^�	$ߠARY�sf"���S@�	�FI��*�$�LINK���!��a_%#�%{q�"XYZ82�*�q�#'OFF���"�"�(%j B�j�4С��n�3FI��%7�q0���j���_J���8%��#�QOP_>$H+5�3�PTB\1�2�C��i�DU�&62�TURN��2r�5`t!}��p��|7FL�`@���m�0�%+*7�^	� 1�. K�	M�&82�Q�2rQ�#�ORQ��G��-( �+p��z�� 3q�E"��T�GOV�@-A��M*�y�4�E:�E@�FW�J��G���D�� o�*� ��A7�P�� y��E�A�GZU:ZU�C�G�ER���	6�E���B�TAFQ��)4�����r'�AX Уa2.q�c�W�c�W �c�W�p�Z�0�Z�0�Z %@�ZK@�Z��Z
!�V � �Y� 
i� i� *i � :i� Ji� Zi� ji�� zi�a�iDEBU{�$v�u��;q�0�"F7O�n�AB���6��CV�z� 
 fr����ukњw�!�w �!�w�1�w�1�w%A�w KA�w��\0��"3LAB"2|EwЄü҂�3 , EE�RVEN� �� $q�_NAǁ!_�PO����` �f�M�_MRA���/ d  T����ERR����~ TYi��RI�V"0�S��'TOQ�T)PL��T��Ѕ_����J � p�PTl X���_V1�b�Q���#��2�2+�����/@�8�p��5�$W��V�j��VN�[�$�@@�� �S���Q�	E�HELL_CFG�N� 5%�Bo_BAS��SRvp\0�K� �S��TJϐ1a�%Α2�U3�4�5�6�e7�8�RO࠘��� � NL:�3AqBn��АACKwv ��)�o�u0iႩ7_PU2�COq��OU��P��ӕ������TP�_KcAR�0��REm��� P����QUE�٩��@���CST?OPI_ALzs���� �TĠ�� SE�M[�w�k�Mw�y�T�Y��SO`��DI����Є�=�װ_T}MK�MANRQζ� E��$KEYSWITCH���Ѱ��HE��BE�AT���EpLE(����&�U��Fd���|��SO_HOM� �O��REF�@PR�i��R� ��C@�O0�p ECO���� _IOCM�4M�k��-��'�O� �D�!ۧH�U��;�M�7��@�3FORC�ߣ�� Q����O}Mq � @EtTxk�U#Po1B�TO�o3B�4x���NPX_AS���; 0ݐADD��(��$SIZߡ$�VAR�TIPRr�q�G�A(ҷ��@
�˨r�t�n�SV��XC����FRIF��R��S%�7�x���N�FѲEАO� x6�PSIڂTEC*�.%CSGL=�T�"�0�&�V�D��>�ST�MT
�o�P\�ByW�@?�SHOWw���P�SV� K�w� ���A00�0 �Q��K���O���_���Ti���5��6��7��8��9��A����@6������20��F�� 
 ����U ����� �����0�� �J@��:�1�G�1T�1a�1n�1�{�1��2��2��2���2��2��2�2��2 �2-�2:�2�G�2T�2a�2n�2�{�2��3��3��3���3��3��3�3��3 �3-�3:�3�G�3T�3a�3n�3�{�3��454��4���4��4��4�4��4 �4-�4:�4�G�4T�4a�4n�4�{�4��555��5���5��5��5�5��5 �5-�5:�5�G�5T�5a�5n�5�{�5��656��6���6��6��6�6��6 �6-�6:�6�G�6T�6a�6n�6�{�6��757��7���7��7��7�7��7 �7-�7:�7�G�7T�7a�7n�7�{�7��M�VP�$�UPD�� � �P���x�YS�LO��� � ���հ�����QTApS�sTƠ��ALU}UL����CU��WFdQ�ID_Lѳ�UHI��ZI�$FILE1_Σ�T�$u�_V;SA��� h��+`?E_BLCK(�8b|g�AhD_CPUQi ��Qi���Sod_R1��ɢR ��
P�W,�d� �aLA��S���c�a�dRUN5��a�d�a�d��5�p�a�d�a�d �T�p�ACC���Xw -$&qLEN~� 3t��&p����Iѱ
�LOW_AXI(�SF1&q�T2mwM��ɢ����I����Q��yTOR.�&p�{DxW��s�LACE����&p�����_MA�uйv�u�w�qTCV�|��wTڱ�;�1�@<ѷt��_��s��J����M��ӠJ����u)���u2q2���������s�pJKцV�K~�か��3ՃJ�0���JJ�JJ��AAL������4�5Xr;�N1�B�N��	��tL�p_�k���"p���{ `5`GROU�P�Y�ӲB$�NFLI�C�ө�REQUI;REv�EBUV�"q���кp2���#pɖx!qxг�� \��/APPRՐC���p�
!�EN�CLOz�,�S_M ���A��u
!q��� 䆣�MC�r;�Xr|�_MGц�C��,`���N��p��BRK��N�OL������Rϰ_CLI��է����JޠѤP��p��p���p;��pD��p6�K���8��n�"q����# ҒMr:ql�Gqz�PATHv��������Rx�������pCNR�CA��է���IN%rUC�pwQ�-Cd�UM�Yop�����QE:p�Gp���~��PAYLOAͧ�J2LHPR_ANqQ�L�`[�W�K�g����R_F2LSHRё�LO\�䱕�����ACRL_@�����޷C�XrH�P�"�$H���FL[EX�!pJ%u� :2Dv�p 4�K�GYq�pPbt|F1Kљխ׃�������E��� �/�A�S�e�w����� y���ф���蘏����$J�ÊT���X���� υ ��څ��[���� 
�� �)��;�D�V��h�z�Y�J��� �� �������QIPA�T��ё��EL4� ��ؘJ���ߐJ�E��CTRޱ��T�N��F�ɗHAN/D_VBp�ѹPn`�� $&�F2���K��ШRSWq?QT�Bj��� $$	M��}�R��E��Uw�H��sA�PH�����Q���A���P��A���Aɫ���j`��D*��DɫP��G�`1)CST��9!��9!N̨DY�`���|�Y� 鰋�KыǦ�J�ч�s�U�ХP��&�/��8�A�J�S�=��� ; �t�.R66N�/QOASYM����Ґ¹���Խ��ٿ_SH�����筈4��+�=�O�JV��h�p'CI����_VI��dHN�u@V_UN!I�ÉD���J҅�B �%�B�̦D�ųD�F�̀���������*Uc�$��Y��H�`�3�XQEN� v�SDIɠS�OwTY��YP��� ��I�1A�Q�äQ�`Bc�S�`�  p�a.a� �[ ME���h�R'R�1TkPPT�0 ) ���Qz�~���0��Xa	iT@� �$DUMMY1���$PS_��RMF��  ��Pf�aLA��YP�jb�S$GLB_T> mU�e�PpQ p���Q�� X	�ɗ`�ST���ߐSBR��M�21_V��8$S/V_ER��OÐ�c��cCL�`�bA5�O�RTPT O�P �o D �`OB���LO˰&uq9c�`�r�0�SYSqA�DR�TP�PTCH>b � ,&��ޥ�W_NA��؀tz�9SR���l =��M�u `�ys�u~�s��s ����������� 0�)�T�"�5�~����B����s�?�?�?D>��XSCRE)�p5�ȐST[�s�}�P!��tX`��r _� Aq� T 	��`ob��a`�l��Ҩ���g�c�O� I�S�c��TX�UE��T� �ñjp^`S<q�RSM_iqmUUNEXCEPlV֑XPS_�a����޳�����޳R�COUx�ҒS� 1�d��UE�tҘR�b9�PoROGM� FL�o$CU�`PO?Q��д�I_�PH�� �� 8џ�_H�EP�����PRY ?��`Ab_�?d�Gb��OUS�� �� @�`v$B�UTT�RV`��C�OLUM��U3�S�ERVx��PAN�E� q��P@G�EU�<�F���q)�$HELPB�l2ETER��)_��m� Am���l���l�0l�00l�0Q�INf��SE@N0�� ǧ1��y��ޠ �)�;LNkr� ��`T�9_B���$H�b TEX�*��ja>�/RELV��DIP>��P�"�M�M3�?,@i�0ðN�jae���USRVIEWq�� <�`�PU�P�NFI� ��FOsCUP��PRI8 �m@`(Q��TRI}Pzqm�UNP��T� f0��mUW�ARNlU��SRT+OL�u���3��O�3ORN3�RA�U�6�TK�vw�V�I͑�U� =$V�PATH��V��CACH�LOG�נ�LIM�B���xxv��HOST�r�!�R��R<�OgBOT�s��IM�� gdSX`} 2����a����a��VCPU_�AVAILeb��EX��!W1N��=�>f`1?e1?e1 n��S��; $BACKLAS��u�n���.p�  fPC�3�@$TOOL�t�$n�_JMPd� �ݽ��U$SS��C6QQVSHIF ��S�P`V��t�ĐG�R+�P�OSU�R�W�PRADI��P�_cb���|�a�Qzr|�LU�A�$OUTPUT_3BMc�J�IM���2p��=@zr��TIL��'SCOL��C���� ҭ�Һ����������o�od5�?��BȦ2Ƣ�0�T��vyDJU2��� �/WAITU����n����%��NE>u�Y�BO� ��� $UPvtfaSB��	TPE/�NEC ��� �ؐ�`0�R6�(�Q��� ش�S	BL�TM[��q��`9p���.p�OP��wMASf�_DO�rdATZpD�J�����Zp�DELAYng�JOذ��q�3 ����v0��vx��,d9pY_���9`7"\���цrP? +��ZABC�u� ���c"�ӛ�
X`��$$C��������!X`��� � V�IRT���/� AB�Sf�u�1 �%�� < QP�/�/
??.? @?R?d?v?�?�?�?�? �?�?�?OO*O<ONO `OrO�O�O�O�O�O�O �O__&_8_J_\_n_ �_�_�_�_�_�_�_�_ o"o4oFoXojo|o�o �o�o�o�o�o�o}� >��AXLMT�s���#  �tIqN&8qtPREO���+vupXuLAR�MRECOV ��)XrzujF }�%�!d������`7�I�[�m�~�,� ��/��uNG5� ��+	 =#�
�ڏ�� PPLIC�5�?�%upՁ�HandlingTool -�� 
V7.70�P/36 ��
�]�_SW2�D�F0<j�W� 43Y�J�|9�K�7DA7?�����
&��a	^-�None��J������ �TG�	�rP_�V�iu�6s��UTO�z"�,tTy.�HGA�PON� %��!.�U���D 1�y� t�x�����y.�K�oQ 1�{  Hp*������	����uq��"�" g�!��Hե�w��HTTHKY��"ٯ����u� ����󿽿Ͽ���� �)�;�M�_�qσϕ� �Ϲ���������%� 7�I�[�m�ߑ��ߵ� ���������!�3�E� W�i�{��������� ������/�A�S�e� w��������������� +=Oas� ������ '9K]o��� �����/#/5/ G/Y/k/}/�/�/�/�/ �/�/�/??1?C?U? g?y?�?�?�?�?�?�? �?	OO-O?OQOcOuO �O�O�O�O�O�O����TOĀ��DO_CLEAND���{S_NM  ɋ����_�_�_�_o��_D?SPDRYR�_��HI!��]@�_}o�o �o�o�o�o�o�op1CU��MAX � bTQNQS�sqXbTB��o�B���PLUGGpb�cWo��PRC4`B�P]klo^�r�O�r=o��SEGF;�K�+�6��_�_}��������ŏ�0�LAPZom�/��+�=�O� a�s���������͟ߟ|�6�TOTAL�v|�y6�USENUZ��g� HXL�NR��R�G_STRING� 13�
�kM,�S�
���_ITEM1��  n󝬯��Я��� ��*�<�N�`�r����������̿޿���I/O SIG�NAL��Tr�yout Mod�e��InpB�S�imulatedޕ�OutT��OVERRW` =� 100��In� cyclHŕ��Prog Abo�r^Õ�>�Sta�tus��	Hea�rtbeat��MH Faul����Aler���� �'�9�K�]�o߁ߓ��� ^S��^Q�� ������,�>�P�b� t��������������(�:���WOR 9���r���L������� ������*<N `r�������PO������ �9K]o��� �����/#/5/�G/Y/k/}/�/DEV� -�/�/�/? ?)?;?M?_?q?�?�? �?�?�?�?�?OO%O>7OPALT��^A ��8O�O�O�O�O�O�O �O__(_:_L_^_p_��_�_�_�_�_LOGRIxp��avO�_*o<o No`oro�o�o�o�o�o �o�o&8J\n�_*�R�ݦqo� �����(�:�L� ^�p���������ʏ܏�� ���PREG bNK��$�r������� ��̟ޟ���&�8� J�\�n���������Ϳ�$ARG_r�D ?	�������  �	$�	[��]���.��S�BN_CONFIOG ��L�K��F�CII_SA_VE  �k��b��TCELLSETUP ���%  OME_I�O��%MOV�_H��¿ȿREP��|��UTOBA�CK��V��FRA:\8�c �8���'`���8�cƅ�'�INI�a@8�^�,�MESSAGz�����|���ODE_D���}�C���O� ��,�P�AUS!��� ((O��J�\� F�|�jߠߎ��߲��� ������B�0�f�t��%�*TSK  �5�c��/�UPDT�����d����XS�CRDCFG 1v��� �������&�8�J�\�n� ��\�n���������� "��F��j|�����/e�2�G�ROUN����U�P_NAܰ��	�2��_ED��1�
��
 �%-BCKEDT-�0�}��pg�ӰQ-2�p8�/�/�8���g2���E/��/��/~/��ED3n/&/�/J/�\.�/"?�/�/ED4 ?�/?�/\.[?�?5?G?ED5�?n?#O�?�\.�?jO�?�?ED6 ZOO�O6O\.�O_}O�OED7�O�Ok_�O�\.G_�_!_3_ED8�_�o�]-�_Vo�_�_ED9Fo�_�o�"o]-�o�oio{oCRoY_Vh�]1��{� LNO_D�ELGE_U�NUSE	LA�L_OUT �V��WD_AB�OR���~�5�IT_R_RTN�ǀH�ONONS)Ю������CAM_PAR�AM 1����
� 8
SONY� XC-56 2�34567890�Y �f�@����?�W�( С���8�h�х�ڎ��HR5ǃ��	���R570�B�Affފ������ڟ� ǟ�"���F�X�3�|����i���į!�CE__RIA_I����5��F��;�Я� ���GP 1]����s�����V�C󠸾�����CO�C ��(���ǀC8��@��H̺�CCX����Ch꺰p��x���� +C�����Ⱥ���+�=�G��ށ��HE>/pONFIG=�f��G_PRI 1�B��tr�����������(�~�CHKoPAUS�� 1���� ,wuj�|�f� �ߊ��߮�������� �.�T�>�x�b���D�O���T���_MORGRP �2?� �\�� 	 �,��P�>� t�b���5�����eҒ.�?a�a�����K(���d�P�V�a�-`�/A�

s��������b&�i��ܦP�DB�����)
�mc:cpmidcbg��:��	�u�	p�U .�n�0� ��d��wC�Ve���g�+/�/f/s/���u/�
DEF ̒�K�)�b buf.txt�/�/���_MC������d,53����|ʇ�Cz  B��p�B��FB�8��B��~C� �Cޢ�D3��u
q�Dzl'D�:�"DrBE�NNEA7E�V�ߓ=F�pg�F=C�F�e,�G���Gp��OG�/�	ބ	6:����4���U(D~���/�ɐʄ3@à1/ � TB�D�V@a � EI�5� F�*� F�G$���F[� GR��kNGl��G����G��&H����G֓�H���߃]��  >�3�3 �ށ� � n^��@߂5Y��Ed��A��=L���<#�
 ��_�*2RSMOFS��.^�9�T1��DE d��,
 Q�;�P�  0_*_>TEKST�"__��R�Q��#o^6C@A�K�Y��Qo2I��BH�0첾@�C�qe�T�pFPROG C%�S�o�gI�q�Ru����dKEY_�TBL  6���y� �	
��� !"#$%&�'()*+,-.�/01��:;<=�>?@ABC� G�HIJKLMNO�PQRSTUVW�XYZ[\]^_�`abcdefg�hijklmno�pqrstuvw�xyz{|}~�����������������������������������������������������������������������������q��͓���������������������������������耇����������������������Eъ`LC�K�l���`�`STA�T�c_AUTO�_DO��O�INDT_ENB;�b��R�QY�K�T2�����STO�~��T{RL�`LETE��ފ_SCREE�N jk_csc 	�Uπ�MMENU 1~i  <�l �ol�K�u���FS�� ��柽�ϟ���R� )�;�a���q���Я�� ���ݯ��N�%�7� ��[�m�������ɿ� ٿ�8��!�n�E�W� }϶ύϟ�������"� ���1�j�A�Sߠ�w� ���߭߿������� T�+�=��a�s���� ��������>��'� M���]�o��������� ����:#p)�+�_MANUAL�ӏ��DBCOu�R�IG�$�DBNU/MLIM�,1e�
�PXWORK 1k�_-�<_N`r�TB_�  m��Y0��_AWAY���1G�@b=�P�_CAL� =���YҀ���`�_�  1!��[ , 

@:&d2/o/�&�Mt��IZP�@P�#ON�TIM��dɼ�&�
�e#MO�TNEND�o$R�ECORD 1'�kU2)?�!�O� ?1-?&k�k?}?�?�? 88�?�???�?c?O*O <O�?�?rO�?�OO�O �O�O�O�O_�O8_�O \_n_�_�__�_%_�_ I_�_o"o4o�_Xo�_ |o�_�o�o�o�oEo�o io�oBTfx�o ��/���� �>�)�7�t�� pu� ����-��͏ۏ��� ��N�`�Ϗ��o���� )�;������8��� \�˟ݟ����;�Q�گ I���m��4�F�X����TOLEREN�C�B�	"�L��Ͱ CS_CFG� ( +x'd�MC:\��L%0?4d.CSVY� �cֿx#A ��CH
�z _/x.�G���},��RC_OU/T )�- z/~��SGN *���"��#�0�3-OCT-25? 11:38���27-MAY���4��]� Z�t�����x.�����pa�m��P�JP��k�VERSION ���V2.0.1�1~+EFLOGI�C 1+� 	d��ٓ��p��PROG_ENB��2��ULS�' ��p�_WRST�JN� ��"�EM�O_OPT_SL� ?	�]�
 ?	R575x#?�74D�6E�7E�50i�d�o�2E�d��|j�"�TO  .�����k�V_� EX�d�% �PAT�H A��A\p��M�_�~+ICT�-F�, '�`ßeg��}�STBF_TTS�(@�	��Eм`���� �MAU��ߧ"MS%W��- )��},t�
��.�!��]l�R �v�����4�SBL_FAUL�y�/��#GPM�SK�ߧ"TDIAb��0����`���!�123456�7890xS�l�P �����//%/ 7/I/[/m//�/�/�/��/�/L0PV ���/�2? X?j?|?�?�?�?�?�? �?�?OO0OBOTOfO�8<x�UMP$�I� �ATR>�Oδ@PME���OY_�TEMP��È��3��4��DUNI�	�w�YN_BRK� 1��x�EMG?DI_STA	���GUNC2_SCR 27[��_�_ �_�_�&�_�_o o2or�nSUQ13y_+?|o@�o�o�olRTd47[�Q��o�o���_ >Pbt���� �����(�:�L� ^�p������� ?Ǐُ �0�,p��+�=�O� a�s���������͟ߟ ���'�9�K�]�o� ��������ɯ���� �#�5�G�Y�k�}��� ����ſ׿����� 1�C�U�g�yϋϝ�ׯ ��������	��-�?� Q�c�u߇ߙ߽߫��� ������)�;�M�_� q��ϧ�������� ��%�7�I�[�m�� �������������� !3EW��{�� �����/ ASew���� ���//+/=/w a/s/�/�/�/�/�/�/ �/??'?9?K?]?o? �?�?�?�?�?�?�?�? OK/5OGOYOkO}O�O �O�O�O�O�O�O__ 1_C_U_g_y_�_�_�_��gETMODE �15'Efa �t|�_GgRR�OR_PROG %�Z%���Hog�TABLE  ��[1O�o�o�o�ZR�RSEV_NUM� �R  ���Q�`a_AUT�O_ENB  �u�SZd_NO�a �6�[�Q�b W *�6p�6p�6p	�6p�`+5pOastHIS�cXa�P{_ALM 17�[� ���6|6`+t���&�8�J�rx_�bp  �[�4q�R���PTCP_VER !�Z�!6oZ�$EXTL�OG_REQ�v9�y�SIZ�܄�TOL  XaD�z�r�=#�
ނ_BWDo�%��f�Q���_DI?� 8'Et�TXa b[�STEPg�y��P���OP_DO�v�$v`FEATUROE 9'EQ��Q�Handl�ingTool �� DER �English �Dictiona�ry�7 (RAA Vis"� Master����
TE0�nalog I/O���p1
0�ut�o Softwa�re Updat�eb� "/�k�ma�tic Back�up
�d
!���ground� EditB�  �25LCa�meraT�FX� w"Lo��ellT���L, P��om�m9�shۡ�h6�00��cou���u�ct��p�pane�� DIF���t�yle sele�ctѡ- /�Co�n��9�onitoir��Hd�tr�?ReliabT�ϣ�(R-Diagnos��Q�	�H��Dual Che�ck Safet�y UIFc�En�hanced Rob Serv���q Hr	ԸU?ser Fr����T_i�xt. oDIO f�fi��u )�\�endܰ�Erru�L��  �prנ*�rO�� �@���ENFCTN Menuİ�v����.fd`�T�P In?�fac�o�  
E�G��p�;�k Excذg��C��High-wSpeܰSki��_  Par+�H��~�mmunic��wons��\ap���urf�?�X�t\h�8U���con�nZ�2Т !�Iwncr��str)��8��M-6�KA�REL Cmd. L��ua��}��~B�Run-Ti�Env�(<�@�I��<�+��s��S/W��"H�Lic�ense���� a�d���ogBook7(Sy>�m)	����"MACRO�s,��/Offs%e\�f����H�!��Y�M1�Mech�Stop ProytZ�3� 5
�{Mi4�Shif\���B6S�Mix�ܰQ����H�Mod�e Switch�Y�Mok���.�� R��Mt�Q�g�� ��5��ulti-Tp������)�Posj��Regi>���  �! �PA�t F�un1��6iB/��R�Num�Y�3��G�P/��� Ad�ju��	�/2HS��)� o(�8�tastu���AD ���RDMޱot�socove&� #e��v�㱗��uest_ 867.��o��\���SNPX b���Y���)�Libr<%�
�rt I����� "����.S�o� ���s in VC�CM����� `j�����㣀/I��� 710�TMILIBX����g��Acc����C/2��TPTX�� �Teln��Y@�����K�PCUne�xceptܰmotn�� ������?\m725�����w�5���  h6�40SP CSX�C�i � j*�� 7RIN��We���g50,��vrlЎزmen" ��fi�P-�a���P��G�rid{�play F O/��? ��fELR;�|�20���ORDK�sci�iw�load�4�1d�st�Patd��CycT�h���oriɰ:�7c D7ata� qu6�2ׁ0�*�������F�RLamc�K�H_MI De��(�����k�PC�φ�Pa�ssword�644��Sp������D#YELLOW �BO�	?1�Arc�%�visu����#t�i�Op�^�! 2ڪ�aO�po�� t���ֶT1o�����H�T��xy�	� �  $�t۠ig���10Ơ 41\�+�JPN ARC?PSU PR+��8b!OL0Sup�2fil� �!��E@�-�;�croc�82p��v���$ 12j�SS0e4�tex�-� I�7�So��t^f�ssag�� e�ēУ�P��,��� "=Tc Virt��v�r��!����dpn��
�J3�SHAD~f0MOVE T�MOS O TԠ�get_va�r fails �l�>PU~1E���� �Hold Bus� %�h��VIS �UPDATE I�RTORCHMA� A�{�vYWELD�TV S ]�DtS:� R741��ou�iPb}�y��BAC�KGROUND �EDIT "RC$R�EPTCD CA�N CRASH FRVR 62z1�SCra��s 2�-D��r ) "���$FNO NO�T RE��RED� �` m ��JO~� QUICKaP�OP FLEN wm41S�Loc���gRTIMQ%�#�F�PLN: FG��p�l m�r`�MD �DEVICE A�SSERT WI�T PCV;PB�A�N#aACCESS� M .pc��Jo��Qui±�KbwldmgUSB$ ���t & rem�ov�� Pg�SMB NUL� ;a|��FIX��C��AC�HIN,QOL�`M�O OPT ՠa>��PPOST0�W�DU C�wQAd�d�`ad���0ioZ�2��$P�`W\0k.$0`O�IN&��P:fix CP�MO-046 i�ssueC�J/aO�-�0�r130Т-� ��vRSET V�ARIABLESx-P{��R3D m��view d��ML��&�ea���b���of FD�5P:~N@x OS-1y0N`�h sc���t���s t�lo��7 W�A�PZ�3 CNT�0 T�/"�Im\R�)�ca �Pu���POT:When�apewB�STY �E�{1t��ptKQd�o GET_�p ��p��VMGR L]Ol�REAd0C~Q W�~1�(�l�s�gD��ECTpLpIN�G IMPR�DR�(p+PB�PROGR�AM�ERIPE:�STARTU� A�IN-;�ӠM/A�SCIIzPÂOF� Lq�DPTTB�: N�pML$m�e P���`:x�mo&�allW`!�ӤTorc�A�U�HC��iLpԸth�`n�@ ch��/GEA��!�tou͐�RC�al��k�Sign�`� ND�ԗThr?esh123��`���09p : MSGs_P�+0er  ��Q�Aܠzeroxn��0 H85�f�RImA�n�2D���rc�0I��OMELa`�pONaP5�  >נSREG:FF-�━ ]�'���KAN�JI��n��J��c��0asn d�!OA �immc �INI�SITALIZAcTI����~1wem����dr+� LB� A�UWqminim�rec[�c!�R����m$�ro -!1>ѮS�ܰir��@�ұJ�1pdETw�� x5`?�I�ow u��~< se 1lc��YbPM���p�Q���R�`vR&�lu\�3�RGe 0�4q�q1#���m <a�arn���ঁBox fyo��*PRWRI�P�W�S��v�09 F��pup�de-rKel2 d�p� j��|`━betwe���IND Q���ig�E snap|�u�s��spo TM�E��TPD#�DO��p#aHANDL �1\k�`vR��ȀD��ny�S�v�Yop?erabil� �TN*�: H � l\pB��Vq�b�R�< p�aj*�c&2O�`FA,��.�-QV7. f.mv��GT�pi��s��� ɠtmL�ine-Rema�rk �� RM-��` W�#SPATH� SA+PLOOS� UIFc�+5f f;ig�pGLA�����Vrp������U�0t�her�V� Trac���tW�\b�s�7��d�t�� n&�@  ���3:����dK�y��it k�8�d�PayR![2y]�ü1: g��]s��dow�XQ��0IS�q�qEMC�HK EXCE yC���MF +��Xah�� 35\k��)���QBt��̐'b���[�c���e� �`k�S�� BU�Gr��cD$`PE!Tp���f�c4��0�XPANSI��D�IG��@OoPme�tTCCRG EN~��CEMENT�A� M̀K {�`H� GUNCHG �`� EXT�P�2�bQS�93 wP8��x�ORYLEAKq  H5gyq�P�LC WRDN �R �O /u�QSPiE=p��G*�V p��$�tn720\3pGRI��A�rT�PMC ETH���pSU7p�`  jy5/n�PENS�P�N,��*P ont��`BROW�`!sR�MV ADDz C�N qDC���PT_3 ALA2@ ����pSVGN EA�RLY�R��ŰH5�7�GaJLAY�ҀE (@M�PP�D�p*@H�S I<`P�OUCH8���rV�F�q�comH�|x ��ERROR� �DE nJ��RO��CURS8pI���N4q�-15y8n7�RSR xP�#aUp���Rqy�T�Fz�;�pk��t�� gՂ�B�S�Y RUNN� � a�`�BRKC�T�!RO�p3@ \3apSТ�AXxP����h8+ q��IS�SUr} sPX�PT�SI�K1M10�_�IPSAFETwY Ck�ECK[� �Á������<#X�� �TWD2�@�@�INV��D Z�Op�5X��t�D�UALy� "M6(�0�"rF#�E��d�PdNDEX F��t*UF�"P�ʀ�0sFRVO1/17 A�PT6�Kt�qFALPTP2+477D6_�P�!;7HIG� CC�t;oSNPX� MM��tq�d~�Vq�q#��
"��DETEC0�Tq*@RRU�qAP�P�5p�9 y�)<9����7T��PdsPp`�2���D�#P��FANUC�p"�I]L02"��U�8�B�	plee�J��hk�3AH�PR�DC"�
�aāp@�@��4A�A�F�b��� �a���I�@���a�G�E<�B�Ccscr�J�@��Ndctrld. �A�N�E�A5��Q���!�`�Df�@�`m�8�78�Q-;�|@�@r�m`�
��PR̠78�@RI�@0q�Q (~\Mp��0t��!>R�@\tQ�	���!�Q�V�St0�3 "	K	`n@���S>V�Rstp�A�@LCF�L���� �Rplcf����J�@�WTamai0�E�@mubov2_mi�@t�O�S�@U`T[tT��AqPr674xSS�hape Gen(���@j�I�[R�`�@b�@T����%q (u�@��II�^�Q�C�a��[�@;Ynrsg0�4�� � 4�Cmr6�@�r5b5�zVnr�etsp "r�P�o�wng0bGCR�E�Ka�ޠ�DA�T�E�k�crea#t.�q�M�a�oks>qgtpad1P��(�tputZj�{�������܆2�@�����Q����sl�o��� �hexH��a�88�ď�keyH��@��pmZb�NR�us�kugc�@UQ�pp�bUZ�dp0aj92�1xSpl.ColAlأcq�\A��RNq̩UA� (J��@ip��_�WA��_�Y��a7�b7�ͦtp[� "TCLS9oKb���clskyh[��s�pkckZd���$��TQ���dA�rx�71�0a- KAREL Use Sp�OFCTN9�a�7l�0s0a�� (���a��@�C�@��q���c8b8"   ��@� Pr	Hr�	   lmatea99�qM��|��E�mcclm5�CLM;�� �j��E�3et���aLM	�h��yasp,���mc_mot�B�N�Ȍ@H����Q��su'��Q��p��䅮���joi#�xߕ��A_log�Z���trc�B����ve�ϓ�v��QWX��~6�finderxS�Center F81�lSw520��hal6rX� (<�r,�Q�Ձfi�Q �r�0�I�ۡ���A�@l��t�q�a "FNDR�Vϳ���etguid�UID�C�@����������a@�nuf;��P���ƞC�B��_z�Ӡo��qG��������l���fndrpTY��2䁴tcp"�,qCP MF�}3Ό@517��6s38 �E��gf6��(���K��Q��-�X��A�t	m6�P�İ��Q���	�͘��t!m�Ĵ�b�@ej���aiex��P@�Aa8�ذ�cprm�A�|�l�_vars� �
��dwc7 TS��/��6��ma�F�Gr�oup| sk E?xchangJ �@��VMASK H5~�0H593 H0a�H5@� 6� 58J�!9�!8\�!4�!�2���"(�/��k���r�� 70a0(�0`�ՁU4U1#SK(�x2�Q�0I�h��)�m�q�bWzR�Dis�playImQ@v�J�@�Q8aJ�!(�P��;� 0a��0���� �@;�qvl? "DQVL�D���qvBXa`�uGHq�O|sC��avrdq�O�xEsim�KЀsJ#st]��uDdX@TRgOyB�BvЀ)�wA~����E�Easy N�ormal Ut�il(in�K�1?1 J553m�0bD2v�Q(lVЀxU)��������k986�#8Uϕ�|�rP "NOR��dw d.a}oKksu�O�W���OY��W`�j0�6�H� me'nuuyP6�M�`wR�X�R577V�90� �RJ989}�4�9b\�`(�fity�����e�<?��&Vsmh`��8�⿠�Sv�q�8���w��pn "MHMN <��ޣx�Ay`�o�3�u �`f�І�x�t��t�RzQ��LV��vP�tm����|I�1{oPx �2�|���I�3I/B�od3stǏًmn���^�}ensu_�L<����h!!��Rt��huserp��0Ҹ�ʐcM�_l�xP�oe�<�рpoper���>�xdetbo/�l> �x���Ps$p�`����OPydspweb ͓��z'R��u�Rr�101&S՟{t�`2�Z4�30�����"�`4�
�4�5��KQp�m[T��dUCalG <�`�Q)p<�}������9;��DA�� �Pr	LATAum�pd�\bbk96M8��68c�fbl�.41969y�9�|�D����bd� "BB�OXêM��sch�ed����m�setauM:�����ff� ��<���n�41�ϒ�<��q�col��|�1�x1c�ؘ���li��X� 0���j��&�8�4 <�{ro5�TP E�l#��ryK42r���;�(T+Q �Rec'�ʈ1Iw�84��x���Ak971���71�;���parecjo��QNS��[T���dXrail| nagek�M ,QjT2 *� (�ĜR%<x�80!bTh��p��4��4�y�Dgl�paxrmr "XRM�g�l��brf{���n��k�l��9turbsp���㧑- �l015	�g�625C�Mh� +���)89��	+��B6��o�ҹ��x��7�q<�����pd? "TSPD�=��tsgl��l�:`dQ���8Bct���K�vrE�aܮ������  1�!���21�`( AAVM �2��0 �@fd T�UP him (�J545 ly)�`8 616 %�VCAM ��CLIO (��0:�5&  (=F\ MSC �Rt"�PBsSTYL��D!28 :2\ N�RE bh SCH�6pDCSU� tpsh �ORSR �rD!0�4�SEIOC�& \fxh 542� LEX"� ES�ETn�8!H ��sh�8 7H �MA�SK�Ø"7>��OKCO*`x�!03"6(�!/400:66$ G6s39.6[8LCH!6oOPLGR703
5OMHCR��0C� h(! �06�A.f8!�54
��00DSWb 588�180 �h!�37 88 (D��"02C24���27 q9�25��2-6��05��9PR�ST bBFR�DMES�!zB�9�30 _ NBA�  6� HLB �3 (~!SM�@ �Con� SPVC� �8!20z��T�CP aram\TMIL A���@PACETPT�X �@p TELON 96��29�%�UECK��r U?FRM et�P!�OR ORP IPL^%CSXC�0j�1�CVVF l F�QHTTP st�A")�I#� CGHP8~ZIGUI�0��hPPGS To�ol� H8�@dj`Z��!@�h!63�%j�@32Q\�31 B��h!96�%R651��Rs�!53 TF�AD�R41�8"1� ��oo�"9��41775�"/@�P�VCTO�@�U�!sh!{80�%PRXY�R��!770 �b8 8�85 ol3P� L� аdi� �`ڳh �LCP{Q� TSS� �b�26:����@C�PE �HT@VRqC~�tQNL ��@002 %��b	0gdis� �`7 <°�a\0�T�`1 �`e=n�b4 652�`)FU02Q0Πo`p2�Ptu�r4 $r�5N��RU0p@ns�e�QJp1 APFiI[ Jp3�g34�g40 alxrE1�t44w46� ts U0  7v�0O��r5�e�p7 p 7"sw�a61:��rY4��r5 QpwGr�`�$�p8R�"sP`tjQ�b�36w77�wL8`�v83���r8�&�:��pOq8�8 "r�key8�9F��a90�91 p�#@���� �D095�g97*pur�A1@d��H�P|P�q1�0QplSqA1p#4��]a!s1@sl༂8�Ӽ�\1�d1�`��v�@{��14p�ae��5 hH2��`�6ޣ��7�f1p@��d�YpCqd�ـ
d�1�`uq��� Cu�1< Oq� ��7ReU	1$ �u1�Pϱ� ���@- WQ158� ase C��9� B��60 82�ń�p���4 (W�ai��`吢!��7�E��8�EU1P`rIo9�<�1��<�2��<�	0��T��l�5HJ�l��cC���9%�GMCR��P�2�`t�Q2@967�QR��8��9Z�2TP�B���P�2P7U5 @�o���
�5�`U���3 w���?A�E$�1��c�qAwl��A��1��512 f���1�u5Р���a5p$��56�+a��Q15h��Ұ�1 @���pp�b[�538 BxaB��|p�4�2�1e1/q5�p�4U5�P16 (߲�Pz��0��8�P�����p�e5`�e5(�/�P`bbf>�X��$Z�U�}5d�\� X¿7 	  ��8� k_kv��79� s�82 &�H�5��E6���p����h ���ñ���3J"�`n��4 3Ȥ59ѧ�6�0t���8��68D0$�$�4 7�����9V�198� ch��ANRS�p��	�C`�90��7�`�|��`�\j670O�`�q�Ӻ�A�C`����q�`���`�t��sg&`�lc���FA`�H��`���`Я���`�hk��`Щ�B`е��o�`���`����`�d�flr��`Ш��� ��o�`���D�;�`�-gEvam����B `г�oќ���`а��>��creexl��ဏ�P��`���|���j�6`�s��prs. `���\���`�7���<���fsgn��P�b�t�at��`�����1B !�svsc�h/  �Servo; S��ule>�7SVS��44�1uӘ_`��� (����ched��,��~���A\�� �� B���B�-AA����cj�� � 5�1`�������p�css "ACS`�&(��6�  �����c el����Q����torcshms�`�- T��Ma`Ѵ���09 �J5;598 JW681s�7� 8 ��b��`Чa����te,s�����/��E�� m��A�RC.�� 1q�4��!� ��C�tc��pA�@t���f� �F����7#�2x�S�E���Utmk �? 60'���RC������� p��96G= '��"H5W����L���\f�� �PATb���`!4U�#!Stmt�E ��� �pMA�!p��8z�2?�in_`Е�(�r�X e/cPA2�`��%����etd�l�vߏ\ovet�o���܏��mmonitr�\��|#F�0st��?.6a�`�PP���! Q8�!y`�`ame �Agrol�c�43��0 �p���01�� 25�  ��`� Pr	H�r	�A�(j818\n; <s�I�B|�2�pMPTP"�|�C�1mocol�� ,��C(�u�'!� �A��̴�8P53��y`Touchs�s�`���!�J5���Ѩ`mP����n[PQ�a,��E�a��IP&
�Pt	h�A`�KF#R�m;�Q�etth�THS�R'�q-�Rt��o "PGIO�#!$s�vISwka�"WK���!�MHqH54J��5w5n/�Sm/���@ 7�*�da��8�`!w/Ac��tsnf Tk�/�#gb�a��(u`��^m�`u�����ܱQp�є�#���HKa<��M��t5Q tZ�a<��dFS5G��4���G�1or��dW��64��tPx���P ����x,��?$����P<�Z4e7�g �"SVGN.ox�copy "CO#�Wj$�O�A�9� "FSG�ѧ�%7��_��5f� wQSWF*!">(�sgatuɀ����_
��tp_TPiDo��9�79�#�dߎ?���h�GAT����!#��  �Гf�` ��"/� �w�Z� �b?6|� ��� �� ���E ���� �chrT� �K6�� ��sms� �o6�ѐ�gtdmen?3 ��&��� ���mkpdt�d2 ���, ���pd�QЕ� ����� ���m?vbkup. �[�xw�С��mkuno���prp���mklh �4��s �niU�<�� �ldvrw���glg�4�� ��棑���aut7�.p б�旐 �ַ������su3� �Ǜ� ��ȷ� ���\ �6�b2 ��?�F��� �����A�4�  ��B ?  946" ��f�� �t\paic\p4k947 ����F#���� �ict3as���pa`���cc:�<��o�����'gen�� � ��F��lnp � ����st1f@��1��wbO�c��Ջ�`��߄�vri �ߢ�а�-T� ��<�p�flow� OP�Ac��ow���R�50qtS �#T� (A��4�#���pѣV�cu3�QF� ��SfI�ac����46�0���s&��pa��!!0���� ���55�b ��o��p���0娿
�aOfcal3�P� ��f��}���`�f��m�	߳�p�d�m�/���a�/��$C`ѷ�� �!? track\P� �0�ine/Rai�l Tr�]TJ�699W�T  (L��8 (`љT.�`�%��D���P0� (��8�4A8��_ɛ�⇒4��P��� �3�b3����alV@ �NT`f���%��Iin]08m���aen���� ��&?5�c@Itst3@��$�� ��`�,R9�%���0��%��popen�ers-OW dD#ev��F�M�6W����|A�Pc"�l!es v� �,��R��V$�Q��0�U<�V$ �k9j ��6��# �����%pwaop/!OPNUp�V ��2celL��8g_��/�6��tscG��$��V!�3z� 5vrop����7`�n(`�V"2 D�a V'O$:S9��� PumpE��jQ��@�r ��!
��@бM SC#�@��)P��AC�`�x�� � Pr����� \mhplu�g�@g�"7P��uXK")㠱io7�CJ0���E�LIO q1�g 7A93շ�5� q9 t����4rb �ST��R��CPJ9s89�P�LSE�'� �e C3Q(P �/Ov���o�P� ?a I1�R���55���f�I1`�tcmio���MIO�����Ut}co1"CL01V� �cBK`io��uM?���Sl�I0�ߢ�DEg �o���f �tI4\onfdtI���ex%�p27�Inte�.TB CoMoo1E��R�(do554# (;r>Ex,��nR##ipc�/>��qp5���
oQé�1��p����7/o���ra�pd�CDV_��r�P�֮��qp2cnd(��s �p��a�o�r@`҄�S��"�c�a�c����2kIԿ?A�p�crt���or0�qd #��"���3p+���D�x�Џ��vr2k�0����AG�.+��c3ho�;�uC��(� �uV630�fwe  P�mී�@���`���TX�� ��d�ch�p "_��(	�3������8����\p3�v����ш�9�3��1 �����lo0w�[ͧ���chk���㳦s��s?Ө0�i�1h���2��i�w����s?1*�-	�:�O��vr������0�'���PFRAPW;at?1rneE�P�sp�& ac5� _A�rbo#�,�a��g@��������Qs<�ICSP+ 9_�x���� ��F��A9PH51IQ93 7��HX6hQ]PVR2`S5��fPR6 iQ�WPR� (P!am S�u�"�A�I>0�tpprg�0����`h�@2atk9�32�!��E�^��asc "8�C��S>i�atp�"�d�@1I��
g�dsblf�ltJA�Qsabl�e Fau�P{C�!��EV0ex/!DSOB (DC��t�$ �p��X 7� �� 5��Q�t3*�~���td9� "!%�(5��sb9኏���\	�6#���@5�p$D@�550-Adju�st PointO"tVJ�Rs�z�䐄���!�X_�Yj��0\sg��4��}7y��\ada�"AD�J���j�Qets{ha<�SHAP�sŭ'jpo�r4�t �!��$ ��C|�	T�k!bRPKAR�/Qiagnost�ì!O!vV66 �J`ew0�(�L���/�&krlde� ��PP���hU b$���r3�Pp?q��ODBG2C��� �@X�o�1U�� ���WT`�@ipJCM��aipper O�pv`1Se}78 (MH GF� ;" :�&##�� a�x�֕$��388C�����#��9.�9C��g##PPk�Q��8�!�_"$ �"��=0%�P��A $���_�#%0AQ�C~2 M�at.Handl�E��!= &�pq MPCLGET�0�1(�3 �Tt&P�Sٰ'�B�1� �B0����&p��H��PP  �'p��@�C7PP	 �TG�tD5�}m�q�Afhnd "F_R?  �����PP	   xT?Q��n�P(Pa��To�P����?�pmpaOx��JP ak925��!2`@O�JRpsQ`B�2�unLHP�Tgse�GSo1�O�W�Q�T��v !�R�Ptpx~���JRdmon.��@��V�!ns�hYvr�QJ�g�Q�o�jY��HS~7sl�f ��pen�PDnR(R&���ɐ823'��ٔq ���g� ���� 1�� St�� ? �c\sltQ �!|QE�P��a�rtPg��P�� �v��"SE�DG8�s0�qtdgY T����vP `ho�s`<`����qc�`g
�e` o�w�a�@o"�ile6�H�e �ȅnR�� �e! j517�>Ճ��J%��e�`��Q!4��Q&�L�!F��J�=�o�5�z/l1�7���_�œ��`C0~C�  ���LANG j��A��������gad���#�jp�.��4�Ē�ib�����Ƒpa���&���?j539.f�,�Ru� EnvA
������3H�z�J9�����h�ФP
Ҕ���2�2����� (KL�n-TimФ�⠤��p��3�TS����\kl>�UTIL"o���~x�r "QMGl���!������1 "���S�T3�\kcmno��SФT2����ut�.�lreadc�}�exY�ܤ�⊸�\��l��Фw�30��2C�*� -�CӀD�E!Ĥ� .��C� �R CV̴�Ҁ�\p��Р���p�tb�ox��.�@�cyc�sL�:�RBTE�v�eriOPTANE���;ӕ�k�e��0��a�ߦ�hg�ߥ��DPN��gp.v�����ptlit���0�4��te\�cy����tm�nu3`�r���5?UPDT��������駣��ite| �� swto�<,���oolB�F"��Y���Q��(q��gr3��䪒��"�䴁Aw������߳��s�������������l<S���bx "O�� ����l����P���A�l\t�� ���ø����	�Col�e!��R C��r���&r �m;`��Cha�ng�Lq�T1 �r�cm3�"��
� 6 ���"����sP7���"L��222���2D457x�� CCFM�|H��accda��Q�c' ��KÕ0���K!����mo!��� ,$Á��!"
��� �/�/����	Y�,$��)�,$sk����m rC%tS1,$+��k1�%unc.,$oñ��1��sub�������1��cce�5/!&@��-/?-W/i&vs� }/�%#�#�/�.C��/� C%
�@? U �&+���F:qt�
pDЃ{ D	  Ux�:7�Dxmov�?81V�@Pe.�P���hPvc5Q�tgeogbdtg_y[tu����P���PxUt�P�Sx�_�^z�_�\var��_�\xy�_�[pc�l`c�P���P�Ue~�Pgripsuao�skuti���ovfinfpo}��o�j�b!�P���Qud\�aX�P�Pc��Rrp�Qnƅ�P�v�P)tm#qƆ�P�v�a+rog�a���Q8�?a+rpal?a{�{spa���P�u�Q�tĊ_xZp�0�osipk�ag3r�ovlcl�ay(�:�t�pT�d �pu?a�c�A����@��KtKa�P����qT�f|rdm��{rin#r���s� �2�ě�|s�Pd�v�tvĈ�v�h�0��ystQn* џ�yt'�1�p���D�p�uϑ#�ul��@o�W6�2�siucpdl�]�o�vr�on��`1L�z�`\�r�΄�il3$|l4��ǉ#q54FyB�Տpg{�`���{wcmס<���wxfer�yY?tlk2pp߿yY�conv��sicn1v�Qʯxag��HώZ�lct`ao�=�p<��׭nit0믁��3������  ��� Pr	H�r	$�	�alϑpm�r&�B�eWa��� f�%������I��� ��u�ͬ�KamT�f�0��c��w��roǁ#� 5�����?� sm�� y�a��y넑������ `����͐ϑ��p��m�Wa�1���A� 6�S�e�X��ψԀQ}� ����������ĥw߉� 西߭���߮�#q0� �rs�ew���1�a��z긱n@�.�۲;��d��ш��  }� �P`	T~$�1 p! P쥰e �e 	tlf@Cь�o/�  ?��%���8�% �x������reg.�C�=��o99 �~@@���$F�EAT_INDE�X  z ���e� I�LECOMP �:���1!�!z$#SET�UP2 ;1%�;"�  N �f!$#_AP2BC�K 1<1) � �)��/�/  %�/�/e4 �/�/ >%�/$?�/H?�/U?~? ?�?1?�?�?g?�?�?  O2O�?VO�?zO�OO �O?O�OcO�O
_�O._ �OR_d_�O�__�_�_ M_�_q_oo�_<o�_ `o�_mo�o%o�oIo�o �oo�o8J�on �o��3�W�{ �"��F��j�|�� ��/�ď֏e������ 0���T��x������ =�ҟa������,��� P�b�񟆯�����K� �o�����:�ɯ^� ����#���G�ܿ� }�ϡ�6�H�׿l���@��ϝ���@)t Px/� 2� *.V1R��߅�*�@�`��F�j�T��PCr�|�߅�FR6:��"��V���z�T � !���K� ��q�SƏ*.Fߢ��	��Ӑ���^����STM ��'����S���iPen�dant PanelS���HI���9����U�������GIF 0;��������JPG��;��]�oR�
ARGN?AME.DTy�E>�\"���R�c	PANEL1Y�%>��e�w��2�A/�//���/�3_/�/� �/p/�/?�4�/I?��7?�/?�?TP�EINS.XML��?>:\�?t?�1C�ustom To�olbar�?Q��PASSWORD�g?w�FRS:\�:O�? %Pas�sword Config{OR��OSO �O�O��_�OB_T_�O x__�_�_=_�_a_�_ �_�_,o�_Po�_Io�o o�o9o�o�ooo�o (:�o^�o�# �G�k���6� �Z�l�������Ə U��y������D�ӏ h���a���-�Q�� �������@�R��v� ���)�;�Я_����� �*���N�ݯr���� ��7�̿޿m�ϑ�&� ��ǿ\�뿀��y϶� E���i���ߟ�4��� X�j��ώ�߲�A�S� ��w����B���f� �ߊ��+���O����� �����>�����t�� ��'�����]����� (��L��p�� 5�Yk �$� Z�~��C �g�/�2/�V/ ���//�/?/�/�/ u/
?�/.?@?�/d?�/ �?�?)?�?M?�?q?�? O�?<O�?5OrOO�O %O�O�O[O�OO_&_ �OJ_�On_�O_�_3_ �_W_�_�_�_"o�_Fo�Xo�_|oo�o�o�`��$FILE_DG�BCK 1<����`��� ( �)
S�UMMARY.DyG�oblMD:�o�*n`Diag� Summary�+8j
CONSLOG qn�=q�ConsoleO log�7kp�MEMCHECKФ�2��qMe�mory Dat�a3�;g� {)>�HADOW(������C�Shad�ow Chang�es���c-��)	FTP������=��qmmen�t TBD;�;g0�<�)ETHERNET0�`n�q~����=qEther�net �pfiguration���B`%�DCSVRF�/��'�@�C�%�� verify� allC��c1p{� �DIFF8�p�0�ůD�%Z�diffǯ{��q��1������J� �X�q�|�	�CH�GD�&�8�ͿD�ܯ�����2Ŀ�����R� `�yτ�GAD�.�@���D�����FY3�ϳ��ώZ� hρߌ�GAD$�6�H���D������UPDAT�ES.$�
�ckFORS:\"�c�>q�Updates �Listc�`{PS�RBWLD.CM���blN��e��pP�S_ROBOWEL\�6o+�=�loa��o ����&���J���n��� ��9��Jo��� "��X�|# �G�k�d�0 �T���/�C/ U/�y//�/�/>/�/ b/�/�/�/-?�/Q?�/ b?�??�?:?�?�?p? O�?)O;O�?_O�?�O O|O�OHO�OlO�O_ �O7_�O[_m_�O�_ _ �_�_V_�_z_o�_o Eo�_io�_zo�o.o�o Ro�o�o�o�oAS �ow�*��` ���+��O��s� �����8�͏ߏn�� ��'��� �]�쏁�� ����F�۟j������ 5�ğY�k�������� B����x�����C��үg�v��$FIL�E_N�PR]����Y�������MDONL�Y 1<��U� 
 ��ۿ(��� L��5���Y��}Ϗ� ϳ�B�����x�ߜ� 1�C���g��ϋ�ߘ� ��P���t�	���?� ��c�u���(���� ^�������$�M��� q� �����6���Z��� ��%��I[����2����VI�SBCK����ų�*.VD�*� OFR:\V� �Vision VD fileV d������� 	/./�R/�v/�// �/;/�/_/q/?�/*? <?�/`?�/�??�?�? I?�?m?OO�?8O�? \O�?�?�O!O�O�O�O �O{O_�O!_F_�Oj_ �O�_�_/_�_S_�_w_��_o~�MR_GR�P 1=��L~eC4  B�`�	 ��lo~li`�۬B��D���fnӺ�MT� ��� ����e`i`a�o�k hb�h�o�dcic.�OL�LX���L�?N��XH�t�E���|�i`@4���B��Az��?�Bf���9�f�l}B+��B+�B,�}B$�!B+���pl}F@� �qhq�y�~g�f�F6�D�Mq�D�� BT��/@���l}?pD�ޒ6���l����5��5���|�l�����ˏ���ڋA�����A��܏e�P���t�  @����@h0?�\	@�B��� ���Ο��+��O� :�_���p�����e;BH` ����	��-�ư��Z��W[C{b/�FX�
�A@���@�3w3@����\��[���ѿ�z��񿋯 �*��N�9�r�]ϖ����<�G�=��<�m]<��+=~�m<c�^��8eN7���7ѷ7��x7;��51�@��	ߤ��?߾d2^`UYb`�b`������F�`Үb` b`�0����C�^o�� �o�o�߸o��o��  ]�(߁�l������ ������#��G�2�k� V�{������������� ��1����- �)������ �0T?xc� ������/') �'/M/_/q/8��/�/ /�/�/�/�/?#?
? G?2?k?V?�?z?�?�? �?�?�?O�?1OOUO @ORO�OvO�O�O�O�O ��_��J����`_*� �_N�_�O�_�_�_�_ oo'oMo8oqo\o�o �o�o�o�o�o�o�o 7"[Fjh� x�t��!��E� 0�B�{�f�����Ï�� �ҏ����A�,�e� ,/���������/�J� ���=�$�a�H�Z� ��������߯ʯ�� �9�$�]�H���l��� ��ɿ��ƿ���#��O �OV� _z�D_V_��z_ �Ϟ_���
�C�.� g�Rߋ�vߛ��߬��� ��	���-��Q�<�N� ��r������� ��)��M�8�q�\��� �������������� 7"[Fk�|� |����֟3� WBg�t��� ��/�///S/>/ w/b/�/�/�/�/�/�/ �/??=?(?:?s?:� LϦ?p��?�Ϧ� O�� $O��T?]OHOZO�O~O �O�O�O�O�O�O_5_  _Y_D_}_h_�_�_�_ �_�_�_�_o��@o
� go*owo�o�o�o�o�o �o	�o-*cN �r������ �)�;�M����� ����ˏݏď��%� �I�4�F��j����� ǟ���֟��!��E� 0�i�T���x���ï�? �?��O��?OO� t�>O������ѿ��ο ��+��O�:�s�^� �ϩϔ��ϸ������  �9�$�6�o�6o��Zo ��R����������5�  �Y�D�}�h���� ���������
�C�U� �y�����d�����:� ����+Q8u `������� ;&_Jo� �����//گ 4/��x�j/4��/X�n/ |��/��/�/!??E? 0?B?{?f?�?�?�?�? �?�?�?OOAO,OeO PO�OtO�O�O���O�O _�O+__O_:___�_ p_�_�_�_�_�_�_o  ooKo6oooZo�oZ� �o�o�o�o��xo
 G2kR���� �����1��.� g�R���v�����ӏ�� �	��-��Q�/*/ ��N/��r/�/ޟ�/� �/)�D�M�8�q�\��� ���������گ��� 7�"�[�F�k���|��� ��ٿĿ���O�O�O�� W�B�{�fϟϊ��Ϯ� ��������A�,�e� P߉�t߆߿ߪ��ߪo ��+�=�a��߅� p�����������  �9�$�]�H���l��� ������������#�G2W}h�p���$FNO �����_�
F0� � } #�1 D|��� RM_CHKT_YP  � �q��� �� ��O=M� _MIN� m�����  �X� SSB_CF�G >� ~�Jl�A�j|�TP_DEF_OW  m����IRCOM�� ��$GENO�VRD_DO�����THR �d�d�_ENB�� �RAVC_GRP 1?3� X�e/��/ �/�/�/�/�/�/�/?  ?=?$?6?s?Z?�?~? �?�?�?�?�?O'OO KO2OoO�OhO�O�O�Op�O�O�O�ROU? �E� q�������8�?�#�O__K_m_o_ꐖ  D3���_Ed�_q�@A��\Bȡ���R��>Y_6 SMT
<#FC-�Ufoxo�o��HOSTC,1�GY?��_ 5	�h�k�o�f�oyeCU gy�z1�������p	anonymous�5�G� Y�k�w��o�o�o��� ���*�<��`� r�������ˏ	��� ��&�8��������� �����ȯگ���M� �4�F�X�j�����ݟ ��Ŀֿ���I�[�m� ρ�fϵ��ϜϮ��� ��}�����,�O�P� ��t߆ߘߪ߼��� /�A�C�(�w�L�^�p� ����ϸ�������� ��a�6�H�Z�l�~��� ��������9�  2DV��z��� ���#��
.@ ������������� ��//g</N/`/ r/�/����/�/�/ ?Qcu��/[?� �?�?�?�?�?)/�?O "O4OFOi?�/�/�O�O�O�O9m�aENT {1H[ P!^O._  `_?_ ._c_&_�_J_�_n_�_ �_�_o�_)o�_Moo qo4o�oXojo�o�o�o �o�o7�om0 �T�x���� �3��W��{�>��� b���Տ��������� A��e�(�:���^������㟦�QUIC�C0�̟ޟ?��1 @��.����2��l��~�߯!ROUT�ER௼�ί/�!�PCJOG0���!192.16?8.0.10	��GNAME !�J!ROBOT����NS_CFG 1�G�I ��Auto-st�arted/4FTP:?�Q?SOB� �?f�xϊϜϮ��?�� �����+�߿�P�b� t߆ߘ�6����� (�J� �1�C�U�g�6� ����������x�	� �-�?�Q�c� ?2?D? ���������) ��M_q����: ���%t��� ��m������� ���!/3/E/W/z {//�/�/�/�/�/6 HZ ?n/S?�w?�? �?�?�?�/�?�?OO <?=O�?aOsO�O�O�O �/
??.?0O_d?9_ K_]_o_�_PO�_�_�_ �_�O�_�_#o5oGoYo ko�O�O�O�O�_�o&_ �o1Cogy ����oT��	� �-�|o�o�o�o��� �o��Ϗ����)� ;�M�_�q���������˟ݟ�ÿT_ER�R I�����P�DUSIZ  j�^���$�>=�?WRD ?޵w���  guest+�}������ůׯ��SCD_�GROUP 2J�� �`�1���!��L_����  ��!�	 i�-	�E����Q�E EATSW�ILIBk�+��S�T 4��@��1��L�FR�S:аTTP_A�UTH 1K�<�!iPenda�n������!�KAREL:*8���	�KC�.��@��VISION SET���u���!�ϣ�������� 	��P�'�9߆�]�o����CTRL L���؃�
��FFF9E3���u���DEFAU�LT��FAN�UC Web S_erver��
�� e�w���j�|��������WR_CON�FIG MY��X����ID�L_CPU_PC����B�x�6��;BH�MIN'��~;�GNR_IO��K���"��NPT_�SIM_DOl��v�TPMODNT�OLl� ��_PR�TY��6��OLN/K 1N�ذ��� 2DVh��M/ASTEk�s�w�}OñO_CFG�Ƙ	UO����CY�CLE���_A�SG 1O��ձ
 j+=Oas �������/�/r�NUMJ�x �J�� IPCH��x��RTRY_C�N�n� ��SCR�N_UPDJ����b$� �� �P��A��/���$J2�3_DSP_EN�~��p�� OBP�ROC�#���	JO�G�1Q� @���d8�?�� +S? /?)3POS�RE?y�KANJI_� Kl��3��#�R�����5�?�5C�L_LF�;"^/�0EYLOGGIN� �q��K1$��$�LANGUAGE� X�6�� ,vA�LG�"S�߀�+����x��i��@�<𬄐'0u8������MC:\�RSCH\00\���S@N_DISP T�t�w�K�I���LOC��-�Dz�U�=#�J�8@BOOK U	L0��`d���d�d��PXY��_�_�_�_�_ nmh%i��	kU�Yr��UhozoLRG_BU�FF 1V��|o2s��o�R���oq� �o�o#,YPb �����������(�U��D/0DC�S Xu] =���"lao����ˏݏ��3n�IO 1Y�	 �/,���� ,�<�N�`�t������� ��̟ޟ���&�8� L�\�n���������ȯ�ܯ�Ee�TM  [d�(�:�L�^� p���������ʿܿ�  ��$�6�H�Z�l�~�p�Ϣύd�SEV� �]�TYP��$���)߄m�1RS�K�!O�c�"FL 1Z�� ����߯����������	�:�TP�5@���A]NG�NAM�$�E��k�UPS PGI|%�1�%}x�_LOAD0�G %Z%CAL_TC� ����MAXUALRM ;'�I(��~���#� QV�#a��CQ[x�@8��n��"�1060\	 �F�	�Ϣ��� ���������� D '9ze���� ����R= va������ ��*//N/9/r/�/ g/�/�/�/�/�/?�/ &??J?\???�?k?�? �?�?�?�?�?�?"O4O OXOCO|O_OqO�O�O �O�O�O_�O0__T_ 7_I_�_u_�_�_�_�_��_o�_,o��D_L?DXDISAc����MEMO_AP�]�E ?��
 �5i�o�o�o�o��o�o�o��ISCw 1]�� �o Td��\no�� �������I� 4�m��f���$����� ����!��E�ƏT� f�:�����ß����� z��ܟA�,�e�w�^� �����~������  �=���L�^�2����� ����߿�r� �Կ9��$�]�o�(t_MST�R ^�͂�SC/D 1_xm�W��� S�������=�(�:� s�^ߗ߂߻ߦ����� ��� �9�$�]�H�� l������������ #��G�2�W�}�h��� ������������
 C.gR�v�� ���	�-Q <u`r���� ��//'/M/8/q/�\/�/�/�/�/�/s�MKCFG `����/��LTARMu_2a��2� �#\`Y>G`M�ETPUT`�"�����NDSP_CMNTs506�5��' b���>�"1��?�4�5POSCFz�7�>PRPM�?��8PSTOL 1�c2}4@p<#�
aA�!aEqOG]OO �O�O�O�O�O_�O�O A_#_5_w_Y_k_�_�_�_�_�Q�1SING_CHK  +O�$MODAQ73d�
?�7:eDEV �	��	MC:>MlHSIZEs0����eTASK �%��%$1234?56789 �o�e�gTRIG 1en�� l��%��?   A$�Üf�YP�a,u��cE�M_INF 1f�>7 `�)AT&FV0�E0N�})�qE�0V1&A3&B�1&D2&S0&�C1S0=�})GATZ�� �H� E��q9m��xAu��� X�������� �� ����v�)���я ��П�������*�� N�����7�I�[�̯ ן���9�&���\� ���g�����i�ڿ�� ����ï4��XϏ�i� ��A���m�������� ��ѿB����ϊߜ� O������ߟߩ���� >�%�b�t�'ߘ�K�]� o߁�����(�_�L� ��p�+����������.�ONITOR�0G� ?ak   	?EXEC1�#U2345T�`789�#��xxx *x6xBxNx@Zxfxrx2U2�2�2�2�U2�2�2�2�U2�33�3�aR_GRP_SOV 1g�y�a(�Q�>�9�?�h����?��<���@�,Ѯ�Hm�a_Di�n�!P�L_NAME �!�5
 �!D�efault P�ersonali�ty (from� FD) �$RR�2� 1h)de�X)dh�
!�1X d�/d/v/�/�/�/ �/�/�/�/??*?<? N?`?r?�?�?�?�?�?�82S/�?O O2ODO@VOhOzO�O�Ob<�? �O�O�O�O_"_4_F_�X_j_|_�_LhR� �1m)9`\b0� �_pb�Q �@D�  �Q?���S�Q?`�QaAI?�Ez  a@o�g;�	l�R	 O0`4b@4c�.a�P�Jd�Jd�K�i�K�J����J��J�4�J~��j0Ea�o-a�@��o�l�[`@�z�b�f�@�S��a�Q�o��c�=�N��
������T;?f�
���m[`��*  �p  ��$p> p�$p���o?��?�����	��o�Bntr�Q�s�kse�}�l�p��  �pu`j7  #p��vks��� 	'� �� �I� �  ���}�:�È6�È=����N��b@�^�d��n�Q���{�RȒx���nN. ��  �'���a�`@a��@�t�@p@hp�n[`CpC0��f0�+pB/pC3}��P�@%��f�oo$|m�/���gA%���. ���z�`�P���QDe���˟��(���m�� �t� O� ru� �4 �xR�c��s� :	e�a�P�` �?�ff  �����7� ��گ쬛af��>搠���iP�P;�e�S�Ea4f�u��>LX��s�b<�	�I<g�<�#�
<2��<D��<��
vo��¯�S��S.����?fff?u�?&�찗d@T���?��`?Uȩ?X����Z���T :z�TB��Wa�з*dů �ρϺϥ���������&�8�#�\�h�+�F . Kߘ�G߼�3���W������G�@ G����X�C�|�g� y���������jZ� ��ￏQ����ߙ� ����3������� /A��t_���
��������F @��@+Fp�IPP�t��%���[`B�0����<z�e�cb!@I��
�M`B@���@`�9@y���?�h� ��@�3�[N���N�N�E���<�/:/L �>���ڟ�A�p��C�F@�S��b/DpX������@�t��%ϑh��`/qG���GknF&��FצpE,�8{�/ F��ZG���F��nE�DE,����/� ���G���F7��F��ED��.��C? .?g?R?d?�?�?�?�? �?�?	O�?O?O*OcO NO�OrO�O�O�O�O�O _�O)__M_8_q_\_ �_�_�_�_�_�_�_o �_7o"o4omoXo�o|o �o�o�o�o�o�o3 WB{f��� ������A�,� Q�w�b���������� Ώ���=�(�a�L�Ѕ�p�����(r!3�3ji��r���ꕢ��3Ա�ڟ�u�4� ����u��P�2�D�&�jb�^�p�1w���������ʯ���ܯ(� �s�P^�PD�c�`�m���y�\������Ӱ�¿Կ���� �.�G����}ϳ� ����홍�U�_�J���$�y.�@�v�d�z� �ߚ�x�4��������� ��D�.�2� �$N[�G�[�^�B�4��B��CH� ^� ���u����������p�h�M�_�q�����������^��^�Y�m�2��
 ����#5GY k}�������h*�� ��>�x}���$MSKCFMAP  ��� �����m�N"ONREoL  6�9�_�"EXCFEN�Bk
7]�FN�C�}JOGOV�LIMkduyd�"KEYk��"RUN���"SFSPDTY�U��v_SIGN|k}T1MOT��z"_CE_G�RP 1n��9\���/���/�/4� �/?�/2?�/'?h?? �?C?�?�?y?�?�?�? O�?@ORO	OvO-OoO �OcO�O�O�O_�O*_�<_#_`_-�"TCO�M_CFG 1oB/���_�_�_
|Q__ARC_�6���UAP_CPL��_�NOCHEC�K ?/ 5�;h9oKo]ooo�o �o�o�o�o�o�o�o�#5GTNO_WAIT_LF'5y"�NT�Qp/��ޙq_ERR�!2q/_�� R_����"�:�L�dT�_MO�sr�}, �{�P_��_�PA�RAM�rs/�������MW��� �=e�345678901.�@�R�)�q� ��_�����˟����ݛLW�3�E�؏i��cUM_RSPA�CE,�������$?ODRDSP�SI&��OFFSET_�CARToݨDI�S�ݢPEN_FILE�I!�Q�v�P�OPTION_I�O���PWORK� t�'�  T�|�C�����6���Z���	 �m���C������RG_DSBOL  ��v����ޡRIENTT5Oj��C���8�=#�?�UT_S/IM_DJ�6	���VàLCT �u�}�����Q��W�_�PEXE���RA�T���� ���UOP ve������������*�8��$���2�#h)deX�)dh�O�X dY�ߑߣߵ��� �������!�3�E�W� i�{������������2n��)�;�M�_�@q�����������<� ����+=Oa�s���X��� O���1m(���(��.�g��"0� �дu�  @oD�  �?���?р��D4 � EzZ3;��	l	 0�ӀS@SM� ��i�i �H)!�H,�H8��Hm�G�	{�G�8��6�MV1��� �C�)����)����Ճ��*  �p  �� > �  �H�/$"�,��B,��Btr�«����¼�/�� �/�"�# �,0 ��� �  z� ߽pj   ���&X�?MU	'�� � 12I�� �  �=��-=���U?g;/�@}?�0~.ѱ��?;Ѳ���H[N	 �?A'M�D�> KC)�f)�" B& ��"O4B+�:�Q��@D1�oo�$����JWAD0�J@�A: �1�E&?��O�O#__G_2]��� �t O�� ru �4 ��R�U��O� :�%S�р~� �?�ff��@[�_�_V_{�o~�b�18р"o0j>�P�Q6YPрZo�WrAd<S�%�>Lw0�#��<	�I<g��<5�<2��<?D��<�׍�l�_�ѳMb�@�?fff?�0?&�p:T@T�q?��`?Uȩ?X�-q�iyBq 5Ya��gI�_ ������!�� E�W�B�{���d������ՏLnpΏ/�ʈG�@ G��U�ȏ y�d�������ӟ���� ���yB=� ��?p� ��/򏸯�߯R�� �'�9��oN�`������~�����ۿƿ�B� ĮD�e�ֿ;�ҿ_�J�?��h�oϨϔ�ϸ��D4��b!�@_@���� ߧ��Ŀ�����%�@I�)�M�`B@��@`��9@y��?���h	� �@��3�[N��N��N�E��<�/�Y�kЖ>������A�p�C?�F@�S���p�X�����@��t��%�h���߉!G��G�knF&�FצpE,8{��� F�ZG����F�nE�?DE,ڏ�������G��F�7��F��ED��Mf��b�M��q� �����������(� �8�^�I���m����� ����������$H 3lW�{��� ���2VA S�w����� �/.//R/=/v/a/ �/�/�/�/�/�/�/? ?<?'?`?K?p?�?�? �?�?�?�?O�?&OO #O\OGO�OkO�O�O�Oz�N(]�3�ji�O�a��	U�E3Ա��O_�a4 ��x%_7_�a�P�Q_�c_ERjb}_�_1w������] �Y�_�_o�_1ol��%P�bPcn~���o��O�o{_�o�oY�`� �o�o,/;M#� f0o�����Y��et�~�i#�1�C�y M�_�����������{b S�Ԏ��	�?�-�c��Mj2���$�VG��z}�B����B��CH�}�9�֟�@����0�B���w�l�~�������Ư�T����\��qQ��U
 ί�0� B�T�f�x����������ҿ���χ��� ���]{x}��$�PARAM_ME�NU ?Յ��  �DEFPULS�E�	WAIT�TMOUTl�R�CV� SH�ELL_WRK.�$CUR_STY�Lj���OPT�����PTB����C���R_DECSN w�Te'�!�3�E�n�i� {ߍ߶߱������������F�A�USE_PROG %P�q%B��V�CCR���UeXÚ�_HOSoT !P�!�����Tt`����������4���_TIMqE�� �T�  A�?GDEBUG��P��V�GINP_FLgMSK]���TR�����PGA�� |��[���CH����TY+PEM�Y�A�;� Qzu����� �
)RM_ q������� /*/%/7/I/r/m//��/�/�/�/�/?��W�ORD ?	���	RS��CP�NS�E��>2JO����BTE���TRACECTL�PvՅZ� a`_ a`{`|�>q6DT QxՅ��0�0D�����0���2��Sc�5{a�0��B���7 �0�2�0B�0B�0젨�2��2�4�4	��4�4�4�4��4�4 ��2�4��4�4�4�4*�4�4�4�4���2�4�4���2!��4"�4#�4���2&
�4'��O&O8OJO \OnO�O�O�O�O�O�OH�O�O�4%X�1(�4U)�4*�4+�4,�4U-�4.�4/�40 _ 2_D_V_h_z_�_�_�_ �_�_�_�_
oo.o@oPRodovb�11�42�4U4�45�46�47�4U9�4:�4;�4<�4U=�4>�4?�4@�4�9�o�o�o�o�o�o �o&8J\n �������� �"�4��1�= �2�D� V�h�z�������¯ԯ ���
��.�@�R�d� v���������п��� ��*�<�N�`�rτ� �ϨϺ��������� &�8�J�\�n߀ߒߤ� �����������"�4� F�X�j�|������ ��������0�B�T� f�x������������� ��,>�bt ������� (:L^p�� ����� //$/ 6/H/Z/l/~/�/�/�/ �/�/�/�/? ?2?D? V?h?z?�?�?�?�?�? �?�?
OO.O@OROdO vO�O�O�O�O�O�O�O __*_<_N_`_r_�_ �_�_�_�_�_�_oo &o8oJo\ono�oV�o �o�o�o�o�o"4 FXj|���� �����0�B�T� f�x���������ҏ� ����,�>�P�b�t� ��������Ο���� �(�:�L�^�p����� ����ʯܯ� ��$� 6�H�Z�l�~������� ƿؿ���� �2�D� V�h�zόϞϰ�������$PGTRACELEN  ���  ��������_UP �y�����������_C�FG z��������<��� �<�Z�l�<�$�DEFSPD {/���a�����IN~'�TRL |/����8Lԃ�IPE�_CONFI+�}>���<�]x�LID(�~/���GRP 1���������@��
=�[���A�?C�C
�XC)��B��r������dL�z�������� 	 �r�N��Ҩ�� ´����B������������A���> �6>7�D_�������� ='�=)���������	 B-��Q�M���  Dz����
��&L7p [�������/�6/!/Z/��
�V7.10bet�a1<�� B�=q�"`ff@���">����!=���͏!A>ff޷!@�ff�"�\�)�"D��?� � �!@�!� �!Ap�#W��h/??*?<?FK;�w����O/ �?K/�?�?�?�?O�? O>O)ObOMO�OqO�O �O�O�O�O_�O(__ L_7_p_[_m_�_�_�_ ��_ o�_$oo!oZo Eo~oio�o�o�o�o�o �o�o DQy{/�#F@ {yw}�y{ ջy�-������ /�Z?l?~?w���t��� ��я��������� O�:�s�^��������� ߟ�ܟ� �9�$�]� H���l�~����_ۯ� �����5� �2�k�V� ��z�����׿¿��� ��1�\n�j�|϶ �������	�4�F� X�j�c�χߙ߄߽� ���������)��&� _�J��n������ �����%��I�4�m� X�����ί�������� ��!E0B{f ������ H�Zό�Vh�ϴϊ ����� �2�D�V� O/�s/^/�/�/�/�/ �/�/�/? ?9?$?6? o?Z?�?~?�?�?�?�? �?O�?5O OYODO}O �O���O�OtO�O�O_ �O1__U_@_R_�_v_ �_�_�_�_�_"4F xBo|����o� �o�o//0/B/;�_ _J�n���� ���%��I�4�F� �j�����Ǐ���֏ �!��E�0�i��O^� ��N�ß՟������ �A�,�e�P�b����� �����o o2oTo.� hozo�o�����o��Ϳ �o
گ'�֯K�6� o�Zϓ�~Ϸ��ϴ��� �����5� �Y�D�V� ��z߳ߞ��������� �1��Uy��:� ���������	���-� �Q�<�u�`�r����� ������T�f� x�n�������� ����7"[F j������ �!//E/0/i/T/f/ �/�/�/�/�/�/?�/ /?A?l�e?w?&?�?�? �?�?�?�?�?OO=O (OaOLO�OpO�O�O�� ��*�O_@RdZ_�l_��$PLID�_KNOW_M � ����A�TSV �v��P�[?�_�_o�O&oo�#o\o�B��SM_G�RP 1��Z� d�I`�oo�$Cf�d����D��TPbj�oLk �f�o"~�U�o> n2T�~��� ��7�4���p�D� ��R���ʏ�������� ��6�
�T��*�����V�QMR�c��mT�EGQK? GR��(� #���[��/�A�S��� ���������$���� W��+�=�O������� ����� ���S�����ST�a1 1�j�����P0� @����E�ϲ��� ������M�0�B�T� fߧߊߜ���������@��7��,�m��2��9���A�<��z�A3�������4���������5)�;�M�_���6x���������A7����������8�(:L��MAD � ���� ��P�ARNUM  ��Ko���SCH
�
 �
��S+UPD��xaq|{��_CMP_�`�� <Pz '�U�E�R_CHK��a��Z���RS���_�Q_MO� �%�_��_RES_G����� ��v/ {/�/�/�/�/�/�/�/ *??N?A?r?e?w?J'��W,g/�?L%��? �?�?N#(��?OON# w�4OSOXON#��sO�O �ON# �O�O�ON#d ��O__N"V 1�x�Uua�@cX��P}p�P$@cW،P}��P@@cV��P��"THR_IN�R���pbA%d�VM�ASS�_ Z�WM�N�_�SMON_QUEUE ��eT��`Ȩ`�N��U�N�V�2`ENqD4a6/NiEXE]o�NeWBE\`>o/cO�PTIO;g?+2`P�ROGRAM %j%1`O_�0b?TASK_I��nOCFG �ox�9pDATAɓ]�B{@ev2w� �����z��+� =�O��s���������^nzINFOɓ��}�!dr��!�3�E�W� i�{�������ß՟� ����/�A�S�e�w�4҇ބ��| �98q~�DIT �B|ׯj~WERFL~h�wS~�RGADJ {�ƪA�  ,��?E�8��Q�IOR�ITY�W���M�PDSP�a�j�U��WvT�OG��_�TG���Rj��TO�E�P1�ƫ (/!AF�PE5 �~��!tcp��>%�!ud�?�!icm<�Q_���XY_<q�Ƭ=�Oq)� *������Op��������� ���<�#�5�r�Yߖ� }ߺ��߳������&�=*�PORT�a��OpA%�_C?ARTREP~`ƭ>aQSKSTA�X!*�SSAV`�ƪ	�2500H80A9u�T毙䕣�ƫ�����`X#�x$�6�m�URGEU`�B��A)WFP�DO�V�2�W�q�?Q��WRUP_DEL�AY �Ưe�RO_HOT�hwR%z�����R_NORM�AL�n��6SE�MI:y�QS�KIP���X%�x 	����� ���X%-;% [mE���� ���!//E/W/i/ //y/�/�/�/�/�/�/ ?�/?A?S?e?+?�? w?�?�?�?�?�?O�?�+O=OOO1U�$RB�TIF��NaRCV�TM�����m@DkCR����A�B
�B}�>�A��@�_�������$������V����HU���o���6��_ <�	�I<g�<�#�
<2��<D��<��
+_ _{_�_)`���_�_�_ �_�_ oo$o6oHoZo lo~oi_�o�o�o�o�o �o�o DV�_z �������
� �.�@�R�=v�a��� ��������׏�*� mN�`�r��������� ̟ޟ�����8�J� 5�n�Y���}���ȯ�� ���A�"�4�F�X�j� |�������Ŀֿ�ӯ ���0�B�-�f�Qϊ� m����������� ,�>�P�b�t߆ߘߪ� �ߧ��������(�:� %�^�A����ϸ��� ���� ��$�6�H�Z� l�~���{�������� ���� 2Vh�� �������
 .@R=O�s �����/�*/ </`/r/�/�/�/�/ �/�/�/??&?28�A�GN_ATC 1���K AT&FV0E02;�ATDP/6�/9/2/9p8�ATA2>,�AT%G1%B9�60k9+++��?,�1H�?,�AI�O_TYPE  �EC/4?RE�FPOS1 1�> K x�O[H/O/�O�MNO`O �O�O�O_�OC_�Og__d_�_K#?_Q_�_ �_�_o�_4o�_Xo�_ Uo�o)o�oMo�oqo�o �o�o�o�oT?x �7�[���� �>��b���!�[� ������{����(�Ï %�^��������A�ʟ e�w���ß$��H�� l����+���Ưa�� �����2�ͯ߯�+� ��w���K�Կo����� ��.�ɿR��v�Ϛ� 5�G�Yϓ�����߳� <���`���]ߖ�1ߺ� U���y��߯����� \�G����?���c� �����"���F���j� ��)�c��������� ��0��-f� %�I�m�� ,P�t�3 ��i��/�:/< O2D2 1�=O� �3/�/�/�/��/�/ ?�/?S?�/w??�? 6?�?Z?l?~?�?OO =O�?aO�?�O O�O�O VO�OzO_�O'_�O�O �O _�_l_�_@_�_d_ �_�_�_#o�_Go�_ko o�o*o<oNo�o�o�o �o1�oU�oR� &�J�n��� ��Q�<�u����4� ��X���󏎏���;� ֏_�����X����� ݟx����%���"�[� ������>�ǯb�t� ����!��E��i�� ��(���ÿ^�翂�� ��/�ʿܿ�(ω�t� ��H���l��ϐ���+� ��O���s�ߗ�2�D� Vߐ�������9��� ]���Z��.��R��� v��������Y�D� }����<���`����� ����C��gM/_$3 1�j/&` ��&�J� G��?�c� ����F/1/j// �/)/�/M/�/�/�/? �/0?�/T?�/??M? �?�?�?m?�?�?O�? OPO�?tOO�O3O�O WOiO{O�O__:_�O ^_�O�___�_S_�_ w_ o�_$o�_�_�_o ~oio�o=o�oao�o�o �o �oD�oh� '9K���
�� .��R��O���#��� G�Џk�􏏏����� N�9�r����1���U� ��🋟���8�ӟ\� ��	��U�����گu� ����"����X��|� ���;�Ŀ_�q����� �	�B�ݿf�ϊ�%� ����[����ߣ�,� ������%߆�qߪ�E� ��i��ߍ���(���L����p���z�4 1��A�S����� /�5�S���w��t��� H���l��������� ��s^�2�V �z��9�] ��.@z�� ��#/�G/�D/}/ /�/</�/`/�/�/�/ �/�/C?.?g??�?&? �?J?�?�?�?	O�?-O �?QO�?�?OJO�O�O �OjO�O�O_�O_M_ �Oq__�_0_�_T_f_ x_�_o�_7o�_[o�_ oo|o�oPo�oto�o �o!�o�o�o{f �:�^���� �A��e� ���$�6� H����Ώ���+�Ə O��L��� ���D�͟ h�񟌟�����K�6� o�
���.���R���� �����5�ЯY���� �R�����׿r����� Ϻ��U��y�ϝ��8��ϧ��5 1� ��nπϺ�8�#�\�b� ��ߤ�?ߡ���u��� ��"��F������?� �����_������� 	�B���f����%��� I�[�m�����,�� P��tq�E� i����� p[�/�S�w �/�6/�Z/�~/ /+/=/w/�/�/�/�/  ?�/D?�/A?z??�? 9?�?]?�?�?�?�?�? @O+OdO�?�O#O�OGO �O�O}O_�O*_�ON_ �O�O_G_�_�_�_g_ �_�_o�_oJo�_no 	o�o-o�oQocouo�o �o4�oX�o| y�M�q��� ����x�c���7� ��[�������>� ُb�����!�3�E�� ��˟���(�ßL�� I������A�ʯe��<����6 1��ϛ� ���e�P�������H� ѿl�οϢ�+�ƿO� �s�� �2�l��ϸ� �ό�߰�9���6�o� 
ߓ�.߷�R���v߈� ����5� �Y���}�� ��<����r����� ��C������<����� ��\�����	��? ��c���"�FX j��)�M� qn�B�f� �/���/m/X/ �/,/�/P/�/t/�/? �/3?�/W?�/{??(? :?t?�?�?�?�?O�? AO�?>OwOO�O6O�O ZO�O~O�O�O�O=_(_ a_�O�_ _�_D_�_�_ z_o�_'o�_Ko�_�_ 
oDo�o�o�odo�o�o �oG�ok� *�N`r��� 1��U��y��v��� J�ӏn��������7 1��ȏڏ� ��}�����ڟu����� ��4�ϟX��|���� ;�M�_��������� B�ݯf��c���7��� [���ϣ���ǿ� b�Mφ�!Ϫ�E���i� ��ߟ�(���L���p� ��/�i��ߵ��߉� ��6���3�l��� +��O���s����� 2��V���z����9� ����o�������@ ������9���Y �}�<�` ���CUg� /�&/�J/�n/	/ k/�/?/�/c/�/�/? �/�/�/	?j?U?�?)? �?M?�?q?�?O�?0O �?TO�?xOO%O7OqO �O�O�O�O_�O>_�O ;_t__�_3_�_W_�_ {_�_�_�_:o%o^o�_ �oo�oAo�o�owo ��o$�oH.�@�8 1�K��oA�� ��o��+��(�a� ��� ���D�͏h�z� ��Ə'��K��o�
� ��.���ɟd�퟈�� ��5�П���.���z� ��N�ׯr�������1� ̯U��y����8�J� \������϶�?�ڿ c���`ϙ�4Ͻ�X��� |�ߠϲ�����_�J� ��ߧ�B���f���� ��%���I���m��� ,�f���������� 3���0�i����(��� L���p�������/ S��w�6�� l���=�� �6���V�z /� /9/�]/��/ /�/@/R/d/�/�/�/ #?�/G?�/k??h?�? <?�?`?�?�?O�?�? �?OgORO�O&O�OJO �OnO�O	_�O-_�OQ_��Ou_[mtMASKW 1�x{oR�_��W�WXNO  ��_�_�^MOTE � �\ita_CFG� �%mpQhuP?L_RANG!aQ�)nPOWER �xu�`1fSM_�DRYPRG �%xz%"_�o�eTA�RT ��n�jU?ME_PRO�o�o�4it_EXEC_�ENB  T-iGSPDpOpWx;dxTDBr�zsRM��xMT_�P�T�`#o�POBO�T_NAME ��Z#�YOB_�ORD_NUM �?�h�QH809  T�O�	�o	O�\�pPO�T� P��a^�	@�M�D|�pP�PPC_TIMoEOUTjo x�PoS232>b1��U��s LTE�ACH PEND�AN��:WYa���� M�aintenance ConsR�ߏV"���KOCL/C�`M�+���L� No Use��+�������NPOf�laYa�/c��CH_�Lp�%nkQ	���MAVAIL�0���h��-e��PACE1 2��[ �Yb�����@S��Yb)�p[ͬ8�?|���� ԯ&�G��\�W����� ����l������ڿ <�M�4��U�Qh͈��� ����0��������@<�M�4�b��o�2t����Ϫϼ�j���� �2���G�h�O�}��3�ߣߵ����߇��� �.�O��d���l�����4����������� �<�Kl/������5������ �7Yh�L������6�� 0�Tv�/�/i/�/�/�/�/��7//)/ ;/M/�/q/�/�?�?�? �?�?�?O��8"?4? F?X?j?O�?�?�O�O��O�O_�O+_��G ;��[ "_��
�P w_oc�_ �_�_�_�_�_onȀG�3mfO@__o_�o��d �`�_�_�o�o�o '9/oAoSnlφHx ��o�o��	��-� ?�Q�Gq�k}�� ҏ����)�;�M� _�q�g���������ѝw `#_ @����po����T�֕ ߟe�w�}�W�X���̯ ޯ�����&�8��� �P���T�f�x���� ���ҿ�F�X�"�,� >�pϲ�tς�
6�����_MODE  y_[�S �_[�Ϭ����O2�[�ĭ���	���ߣ�CW�ORK_AD-�	�,߸��R  �_[O@D���.�_I�NTVAL-�tD��8�R_OPTIO�Ne� 8��$�SCAN_TIM�,���8���R ��(�30(�L�8��P�R���� ����A���������e�σ#�2�Q�����d]�T�d����㵛@��������h�Wx���P�U���@OA,> D��Ohz�� �����
���B��(as�pK���A;��o�T��Ap3�?t��Di����>��  � l#�~E ������//+/=/O/ a/s/�/�/�/�/�/�/ �/??'?9?K?]?o? �?�7��?�?�?�?�? �?O!O3OEOWOiO{O �O�O�O�O�O�O�O_ _/_�?�?0p_�_�_ �_�_�_�_�_ oo$o 6oHoZolo~o�o�o�o��o�o�o�e  0 �RW�=Oas� �������� '�9�K�]�o������� ��F_ۏ����#�5� G�Y�k�}�������ş ן�����1�C�U� g�Ə؏f_����Я� ����*�<�N�`�r� ��������̿޿��0�&� w,  WZ� l�~ϐϢϴϾ����� ����+�=�O�a�s���ߗߩ߻����� ���O���0�B�T� f�x����������a�������H�� �G�	12345678K�_���Q �������������	�&8J\ n�������� �"4FXj| �������/ /0/B/T/f/x/�/� �/�/�/�/�/??,? >?P?b?�/�?�?�?�? �?�?�?OO(O:OLO {?pO�O�O�O�O�O�O �O __$_6_eOZ_l_ ~_�_�_�_�_�_�_�_ o=_2oDoVohozo�o��o�o�o�o�o�oP� I�+s0oUgy���Cz  Bp���   ���2��z�$SCR_�GRP 1�(��e@(�l����@ >0� +�9��	  �s���DqF�B�)��O� �M�;�t���-�	�C������E�����q�ǌLR� Mate 20o0iC _�90W���W�LR2C �`�V��V�V��
6�l�E��%�R�0�ǃF�q��E�S�	�D�������ҟ���.�����/�$�7� q�Z�l�?��6����C�ԯ�xƯ�vh:�,>�BǛp� ��7�r�A�pF�  @��^��@��n�  ?�����H�p��I��F@ F�`�� ɿ���ؿ���!�G� 2�k�VϏ��^�����0�Ϸ�����B���~� /��S�>�w�b�t߭� ���߼�����﨎�@
�]��L�^�_�
h���|ㆱ@��=��a"��@�r���B� �[�90��w�p�EL_DEFAU�LT  ����|�.�M�IPOWERFL�  &�F�-�S�W7FDO;� F��q�ERVENT 1O����D�p�L!DUM_E�IP�����j!?AF_INE:����z�!FT�����1!!�V �� }!RPC_OMAIN~`�l���VIS�_	���!TPP�U��da!
�PMON_PROXYb��eP�(�{��f��!R?DM_SRV���9g�E/!R"�e/���h4/�/!
� M����i�/�/!R�LSYNC�/9�8�/)?!ROS��P<�4?u?D�? #f?x?�?�?�?O�? /O�?SOOwO>OPObO �O�O�O�O__�O=_�_a_(_�_��ICE�_KL ?%��� (%SVCPRG1�_�Z�U�s�_"�]3�_�_�P4"o'o"�P5JoOo�P6rowo�P7�o�o�P��ol	9�o�k�T\/�Q �_?�Q�_g�Qo� �Q<o��Qdo��Q�o ��Q�o/��Q�oW��Q ��Q-���QUϏ �Q}���Q���Q� G��Q�o��Q����Q E����Qm���Q��� a���_�R�P�_�PZ� ���q��ǯ���֯� ��3��W�i�T���x� ����տ������/� �S�>�w�bϛφϿ� �ϼ�������=�(� a�L�sߗ߂߻ߦ��� �����'�9�$�]�H� ��l�������������#��Z_DEV ����MC�:+�|h=�O�UT/6�N�9�REC 1�|�6���� 6� 	 u6���  
6�����b��������������.b��
 �Z�6 s��A��{���'��6�)J6�{6�Uz6�BO�������O����{�|�R �V r�Z� �  x���M % �� �6�6�[�a6�T&��XO� �6��?� �N����*������ mQP�v 6�6��=6�[6��T���TO� �6��*� u�3/��òVH���һ ?�  �"/�*=�6�z6��~/��e�� �6�6� z�/�/F/~KV��(6�t6�6�u�ю6�5��Z*? �6�kO��C6�b6�qR?�?�/~NV�9	���z?6�P6�>�:	�?d:D6�6�oX�?7O�?��V"6�Ui��b6�����&O��6�6�/�6�|N? O�QQE*O�پ �6�$� )F(.O@ORH�V*���4�!0�@��O����H�6�_._6�CJO�о ��O�V_�_�O��Q倍%0��~_@Z<(NT�g[�vT$o;o��_�&6�M�V����W6�*o�s"�6�6�RNT[��o�; �b1O�" �o�o�>�O �m�i* N<r`��� �����&��J� \�>���n��������� ȏ�����4�"�X�F� |�j�������֟ğ�� �
�0��T�6�H��� x�����ү������ ,��<�>�P���t��� �����ο��(�� 8�^�@ς�pϒϸϦ� ���� ����6�$�Z��H�~�lߎߴߌ�V C1����0�o�����   -����h�1�_TY�PEx�;�HELL_CFG �J�6��� ���RS�a������ ����:�%�^�I��� m���������� V!��0���%! Oa�6�8�1u1!Al�u1u0��g7!Qd�ygV�HK 1�d� �" 4]Xj|��� ����/5/0/B/�T/1�Y�OMM �d�/U�FTOV�_ENPD���M�O�W_REG_UI��/T�IMWAITp�"}`�+OUT�&����)TIM�%;��0?VAL?�#_UNIT�#g6M��MON_ALIA�S ?e�) ( he�Ѿ?�?�?�? O�f�?3OEOWOiOO �O�O�O�O�O�O�O_ _/_A_�Oe_w_�_�_ �_X_�_�_�_o�_o =oOoaosoo�o�o�o �o�o�o'9K �oo����b� ����5�G�Y�k� }�(�����ŏ׏鏔� ��1�C�U� �y��� ����Z������	�� Ɵ?�Q�c�u���2��� ��ϯ�󯞯�)�;� M�_�
���������d� ݿ���%�пI�[� m�ϑ�<ϵ������� �Ϩ�!�3�E�W��h� �ߟ߱���n������ �/���S�e�w��� F�����������+� =�O�a���������� ��x���'9�� ]o���P�� ���5GYk ������� //1/C/�g/y/�/ �/�/Z/�/�/�/	?�/ -???Q?c?u? ?�?�?�?�?�?�3�$SM�ON_DEFPR�O ����
A �*SYSTEM*�  �l��4R�ECALL ?}�
I ( �}6�copy frs�:orderfi�l.dat vi�rt:\temp�\=>asusv�ivobook1�4:7704 4�  0 7818�5 �A�O�O�O  ;}.JF*.d^OpN�yO�O_._�E
xy�zrate 61 �O�O�O_�_�_�EJWc_}Qj_|_�_o�1o�B9JDh:\s�upport\*�.*WTTi=>27�983872:301555o�o�o�M8JBXSoutp�ut\calpo�int.pc md: overqo�o%�N5�otcp_1�owj ���HZs2as���(��K7��`_\p.ls��h������M�!ersrch �0x160002o� l�~��!�3�F��X�j���������BAJBg�\�tpN�֔k���s���0�CkQO[Qmpbackb_�R�(�����L0ʔb�@^e�f�uI{����0��C4xJ�:[hݥ\`��Q@���������pJ�aR� d�v����$Ϸ�I�[� ���`ϓϥϸ�ʟN� � ��#�5��Z��5  ߑߣߵ�H�Z� ����!�3�Ư��� �����D�׿�z� ���/�¿������
� ����@�R�d�zg�� #5����c�~�� �F�aj�|�1 ��W�i�����B� Sex��/-/���� ����/�/�/�o�o�o �m�/?'?:/L/^/� ?�?�?8?J?�n?�? O#O5O�?Z?�?�?�O �O�OFX���O_ 1_��O�O�_�_�_ BS_�x�_o-o� ��_�o�o�o>OPO bOt/�o)�O�OW_ no��:_L_gp_���%�6��$SN�PX_ASG 1߶���U��� P��'�%R[1]@g1.16���?���%������Џ��ŏ� ��<��`�C�U��� y���̟���ӟ�&� 	�0�\�?���c�u��� �����ϯ���F� )�P�|�_�������ֿ �����0��%�f� I�pϜ���ϣϵ��� �� �,��P�3�E߆� iߐ߼ߟ�������� �� �L�/�p�S�e�� ������ �����6� �@�l�O���s����� �������� V 9`�o���� ���@#5v Y������/ �/<//`/C/U/�/ y/�/�/�/�/�/�/&? 	?0?\???�?c?u?�? �?�?�?�?O�?OFO )OPO|O_O�O�O�O�O �O�O_�O0__%_f_ I_p_�__�_�_�_�_ �_ o,ooPo3oEo�o io�o�o�o�o�o�o��o L/tH�PAR�AM �U��_� �	�PzP��t�p@�OFT�_KB_CFG � �s[��tPIN_SIM  U���v����pH�R�VQSTP_DS�B�~�rM��xfpS�R ��{� &�  AL_TC�u���t�vTOP�_ON_ERR � �t�y��PT�N �u��A��RINGo_PRM�� fp�VDT_GRP �1�uyɀ  	 �w�x2�D�V�h�z��� ����ԟ����
�� .�@�R�d�v������� ��Я�����*�<� N�`�����������̿ ޿���&�M�J�\� nπϒϤ϶������� ��"�4�F�X�j�|� �ߠ߲���������� �0�B�T�f�x��� ������������,� >�e�b�t��������� ������+(:L ^p������ � $6HZl ~������� / /2/D/V/}/z/�/ �/�/�/�/�/�/
?? C?@?R?d?v?�?�?�?��?�?�?	OO�sVP�RG_COUNTƷv���u4BEN�B��/EMYC�tfO_�UPD 1��{8  
O�r�O�O �O�O�O
__E_@_R_ d_�_�_�_�_�_�_�_ �_oo*o<oeo`oro �o�o�o�o�o�o�o =8J\��� �������"� 4�]�X�j�|������� ď�����5�0�B� T�}�x�����ş��,EYSDEBUG>@ʣ@�Аd�I�SP�_PASS>EB�?�LOG �V�E�CА͘�ڟ  ��AБ
�MC:\0���1�_MPC6��E��į�A�m�� �A��SA/V �9�V�q��Еx�SV�T�EM_TIME �1��K (  [�Гy͘%���T1SVGUNS��@?E'�E���A�SK_OPTIO�N>@�E�A�A��BCCFG ��K�� ���` �J�B�-�?�x�c� �χ��ϫ������� �>�)�b�M߆�qߪ� �ߧ��������(�� L�7�p��Еn�� o�����]����<� '�`�鮀���U����� ����������* ,>tb���� ���:(^ L�p����� ���/ /2/D/�h/ V/x/�/�/�/�/�/�/ 
?�/.??R?@?b?d? v?�?�?�?�?�?�?O O(ONO<OrO`O�O�O �O�O�O�O�O__8_ �P_b_�_�_�_"_�_ �_�_�_�_"o4oFoo joXo�o|o�o�o�o�o �o�o0TBx f������� ��*�,�>�t�b��� N_��������(� �8�^�L�������t� ʟ���ܟ� �"�$� 6�l�Z���~�����د Ư����2� �V�D� z�h�������Կ¿�� ���"�@�R�d�⿈� vϘϾϬ�������� *��N�<�r�`߂߄� ���ߺ�������8� &�H�n�\����� ����������4�"�X� �p���������B��� ����BTf4 �x������ �,P>tb� ������// :/(/J/L/^/�/�/�/ n��/�/ ??$?�/H? 6?X?~?l?�?�?�?�? �?�?O�?2O OBODO VO�OzO�O�O�O�O�O �O_.__R_@_v_d_ �_�_�_�_�_�_�_o �/0oBo`oro�oo�o��o�o�o�o�f p��$TBCSG_G�RP 2��e�  � q� 
 ?�   K]G�k���@����$r+s�2|�d0 �@�?� q	 HBH�L���\��B   �CQ�w���P���o�D��΍A���H����A��T�q	�Ԋ6f)f��6�@ pC��^�c@�6�|��C�^� `�~���u������v�� �'���R�o�:�L�x����ƫ?Y������	V3.0�0Cr	lr2cƣ	*���r�\Цő�33 p4�Ɯ� H��I�  �^�����$qJCFoG ��e<qY ?p�����r�9������ ��`�A�,�e�Pω� tϭϘ��ϼ������ +��O�:�s�^߃ߩ� ���߸������ �9� $�6�o�Z��~���� Cr]`�������+�� ;�a�L���p������� ������'K6 [� q��o�� � �$H6l Z|������ /�/ /2/h/V/�/ z/�/�/�/�/�/
?�/ .??R?d?Zo|?�?8? �?�?�?�?�?OO<O *OLOrO�O�OTO�O�O �O�O�O_&_8_J__ n_\_�_�_�_�_�_�_ �_o�_4o"oXoFoho �o|o�o�o�o�o�o�o 
TBxf� ������?� � 2��b�P�r�t����� ����Ώ��(�:��� ^�L���p�����ʟܟ ���� �6�$�Z�H� ~�l�������دƯ�� � ��D�2�T�z�h� ����¿���Կ���� 
�@�.�d�RψϚ�D� ���ςπ����*�� N�<�^�`�rߨߺ��� �������&��J�\� n��:�������� ����"��F�4�j�X� z�|����������� ��0@fT�x �������, ��DVh��� ����//:/L/ ^/p/./�/�/�/�/�/ �/ ??�/�/H?6?l? Z?�?~?�?�?�?�?�? O�?2O OVODOfOhO zO�O�O�O�O�O�O_ 
_,_R_@_v_d_�_�_ �_�_z�_�_��_<o *o`oNo�oro�o�o�o �o�o�o�o8&\ J����p�� ���4�"�X�F�|� j�������֏ď��� ��B�0�R�T�f��� �������ҟ���� >�,�b��_o����H� v���ί��(��L� :�p�������d�ʿ�� ڿܿ�$�6�H�Z�� ~�lϢϐ��ϴ����� �� ��D�2�h�Vߌ� zߜ��߰�����
��� .��>�@�R��v�� �����������0� B���r�`��������� ������&8J�n\����  9� � �����$TBJOP_GRP 2Ũ��  G?���{� 0'�Z@�U � �:p�� c+	 �BL  �?Cр D�+���?fff�:�lB ��f�f@��33D  ��/'��@/R,cd%9<�}b�Y��?�z ����/�AЮ'D� $�3/��%�/>�*9�P�A�y}@����C�* x0�/-?A6ff@5�0!D/cR(�� d2]?o>p!�9%1� �1�?�?@	1�4L?R$�&��1�?S#333|B,8���?� c?Lv00+B�2C�;OMO�?�?�*�O >��ff�AB�� $O6O�O6/�E�O7_ �O_6_g_B_�O�_�_ �_�_�_�_�_�_o0o`o(oVo�o�C����ahe	V3.�00flr2ce*�`e��o�g� E���E��A E��E���3E�iNE��!hE�فE�ۑ�E�I�E���E���E��rF�F��FM(F��5FBF�aOF�\F�"f�bz  E��@ E�� E��� E�  E}�^p�� E�Zp_�� E�Vp�^p��Vp� F  � F� F$� Fj` F�@� F�P F�`� 9�IR9�%opl�uj��
�r��s�A?!��ESTPARS��p�%	HR;�A�BLE 1�$��&��w T��y
&�&�&���&�	&�
&�&�u��&�&�&��qU�'RDI]�$t��� ������΅6�O>�P�@Z�l�~�����V�S<�"  �c�u������� ��ϯ����)�;� M�_�q���������� ;�?�n�������� ŏ׏�����V�ಿNUM  �U$l�  �p��pV�_CFG ����v�c@IM?EBF_TTA�q�8"N��VER�s�z!��R 1�O
 8�o�� 2~� � �  f�x� �ߜ߮���������� �,�>�P�b�t��� ��������)���,�H:�L�K�_��8�@"��
MI_CHA�N� "� ��DB'GLV! �"����ETHERADW ?� �#��^�\�$��RO�UT5�!!�VtGSNMAS�K "255�.��c��OOLOFS_DIA������ORQCTRL �C���>8-bt��� ����//U�R�$/6/k/7�PE_D�ETAI��PON_SVOFF��}#P_MON ���� �2w)STRTCHK ��=~"VTCOM�PAT�(|$� FPROG %�%  AL_TC�P?r.�PLAY�B��*_INST_�M�  �<Y'�4UqS5�-??2LCK�<��;QUICKMEx���??2SCRE@�
tps��`?2�11@6I��G@_�KI\�*9��SR_G�RP 1� �k�ҶO�J��O�O�O_�O/_^� �V_dZ)Qq?�_y_�_ �Uho�_�_�_�_#oo Go5oWoYoko�o�o�o��o�o�o�oC	�1234567�8Wi6�X0E1���K
 �}ip�nl/�pgen.htm�_��� ���(�Panel setup�}?V�h�z������� E�;������ 0�B���f�ݏ������ ��ҟ�[�m��,�>� P�b�t������ί ������:���^� p���������/�A��  ��$�6�HϿ��� �Ϣϴ�������a�� ��2�D�V�h�zߌ�߾t>UALRM�0G� ?
   ��������"��F�9� j�]�o��������������SEV  ���>���ECFG ��-��eQ}An�   B�y4
 �y3���� ��������1C�UcJ�B��+ P��_��IC6?M;W (% ��� � =(aL�p������/��4 ���/I_@H�IST 1��) � ( ; ���%/SOFTP�ART/GENL�INK?curr�ent=edit�page,,1 �`1� �/�/�/�/�*�y(�/�%menu�"955� �/E?W?i?��/
??148,2 _XY4?�?�?�?X?�?�=53�!Z�?@OOaOsOOO�?0>O �O�O�O_�@'�O>34� � 4�OX_j_�|_�L,_�.CAL �/�_�_�_o_)_� 71� MV�_^opo�o�m���!��o�o �o�o�C�oCU gy��,��� �	���?�Q�c�u� ����(�:�Ϗ��� �)���M�_�q����� ��6�˟ݟ���%� ��Ɵ[�m�������� �oٯ����!�3�E� H�i�{�������ÿR� �����/�A�пe� wωϛϭϿ���`��� ��+�=�O���s߅� �ߩ߻���\����� '�9�K�]��߁��� ������Ư���#�5� G�Y�k�n�������� ����x�1CU g�������� ��-?Qcu ������� /)/;/M/_/q/�// �/�/�/�/�/?��/ 7?I?[?m??�?�/�? �?�?�?�?O�?3OEO WOiO{O�OO.O�O�O �O�O__�OA_S_e_ w_�_�_*_�_�_�_�_ oo�_�_Ooaoso�o �o�o8o�o�o�o�':�$UI_P�ANEDATA �1����Wq�  	��}  frh/c�gtp/widedev.stm3������|)  ri~�0hp�(� :�L�^�p�������� ʏ��� ��$��H� Z�A�~�e�������؟~6� � �� # Q�� �'�9�K�]�o��� ���ɯۯ����x� 5�G�.�k�R������� ſ��������C�U�<�y����Ys�� ����������f�7� ��[�m�ߑߣߵ�� ���������3�E�,� i�P��t������� �����Ϣ�S�e�w� ������ ���D��� +=Oa���l ������' 9 ]D��z� *�<���/#/5/G/ �k/}/���/�/�/�/ �/�/b/??C?U?<? y?`?�?�?�?�?�?�? 	O�?-OOQO���/ �O�O�O�O�O�OFO_ �/;_M___q_�_�_�O �_�_�_�_�_o%oo Io0omoTo�o�o�o�o �o�o�opO�O3EW i{��o�$_�� ���/�A��e�L� ��p��������ʏ� � �=�$�a�s�Z��� 
͟ߟ���'� z�K�]���������� ɯۯB����#�5�� Y�@�}���v�����׿��п���1Ϥ���}�B�{ύϟϱ�����)i���m���&�8�J� \�n߀��Ϥߋ��߯� ������"�	�F�X�?� |�c������i�������$UI_PA�NELINK 1����  ��  ���}1234567890/�A�S�e�w� ����i�-��������� ��7I[m��)	)���p��+�  SOFTPART/GEN��?CONFIG=�SINGLE&P�RIM=mainedit �+�=)
��M=wi?ntpe,1� ��X��//*/ </��r/�/�/�/�/ �/d/�/??&?8?J? �/X?�?�?�?�?�?`? r?�?O"O4OFOXO�?�fO�O�O�O�O�O�� 0,  	 E�or��#^Pco 
_K_.Wg_y_\_�_�_ �_�_�_�_	o�_-o?o "oco��vo�o�m*� ���o�o+=0 �ogy����P ��	��-�?���� đ]�i���������� Ϗ��b��/�A� S�e�w��������џ ������+�=�O�a� s��������ͯ߯� ���'�9�K�]�o��� �����ɿۿ����� #�5�G�Y�k�}Ϗ��G �Ͻ�Lo��������� ;�M�0�q߃�fߧߊ� ��������dq�q� �oM��o������� �����&�8�J�\� ��������������� [�m��4FXj| �ϲ���� �BTfx�� +����//� >/P/b/t/�/�/�/9/ �/�/�/??(?�/L? ^?p?�?�?�?5?�?�? �? OO$O6O��ZO�� ~O�OsO�O�O�O�O�O _ __D_V_9_z_]_ �_�_��_C��_g�o .o@oRodovo�o{��o �o�o�o�o�o*< N`r����? ����&�8��?\� n���������E�ڏ� ���"�4�F�Տj�|� ������ğS����� �0�B�џf�x����� ����үa�����,� >�P�߯t��������� ο=O�ϓ_(�:�� ^�Aςϔ�wϸ��ϭ� �����$��H�Z��_ {��_��o�������� � �D�V�h�z�� ���?�������
�� .����v������� ������q�*< N`������� �m&8J\ n������� {/"/4/F/X/j/� �/�/�/�/�/�/�/�/ ?0?B?T?f?x?翜? �?=��?�?�?O�?,O >O!ObOEO�O�O{O�O �O�O�O�?[�]���K]��$UI_POSTYPE  e�� 	;R�K_O__QUICKMEN  l[�:_�_^QRESTO�RE 1�e��  � ���Boo8im3o\o no�o�o�oGo�o�o�o �o�o4FXj| 'o������ �0��T�f�x����� ��Q�ҏ������ '�9�K����������� Οq����(�:�ݟ ^�p�������Q�[�ů ׯI���$�6�H�Z�l� �������ƿؿ{��� � �2�D��Q�c�u� 翰��������ϛ�� .�@�R�d�v�ߚ߬�������XWSCRE��P?�]uw1sc�Pu2�U3�4�5�6��7�8�]RUSE�R����T���k�s'��4��5��6ʆ�7��8��]PND�O_CFG ضl[  �P ]PP�DATE h���None �V]PSEUFRA_ME  �D�����RTOL_AB�RT�[R�ENB�(��GRP 1���Y�QCz  A�~�|��A|������������������PU�H���7�MSK  �K�S7�N�%�1UT%�ߌZRVI�SCAND_MA�XII�3�� FAIL_IMGI �6P��@#S�� IM�REGNUMI
���SIZI�P����,�ONT�MOU'�K����&���c�� �V�s�FR:�\� � �MC:\(\LO�GhB@�� !�{�����Ez? MCV��oUD1 &EX	+��C6PGe��lYz�0(yQ=���c/���`/r/�/�/�/ �/�/�/�/??&?8?�J?\?�PO64_r���pVn6�5�!�LI��:�8�1V��<f@�7�?�w =	�8SZV�>w����7WAI�?��STAT ܄k��@@��O�O�J$��O�O� �2DWP�  ��P G��@tR1�H�O�_�JMPERR 1��l[
  ��23�45678901 RV��v_i_�_�_�_�_ �_�_�_oo<o/oAoxro�$ MLOWQN8�� �_TI/���'� MPHASOE  �����`��SHIFT%1=N+
 <plz 2�e7pGY� }�����$�� �Z�1�C���g�y��� ؏��������D����e���k�	VS�FT1s3V� MN�� �5A�� p����A�  B8*�������pǓ��b�����5 h�ME�@�K��i��1QN&%���aM���N+�@��	 �$N@TDINGEND34J�OH +h�1~�S��e��`.I����GO�߭ q����⪰��ϯc�RELE�aI�G�.�@J�_ACTIV�TƲ��A �`mS����ƲRD�0�����YBOX ����dϻF��@2�~��190�.0.��83n����254n��a���x0~������A�robot���o�   px�7߻Epc�� X�Kئ�F���H۠���^��ZABCd��k�,KP���BV����.� �'�9�K��o��� �����������<���	Z�Aǜ�