��  ë�A��*SYST�EM*��V7.7�077 2/6�/2013 A�Q  �����ABSPOS_G�RP_T   � $PARA�M  	�  �ALRM_�RECOV1   $ALMO�ENB��]ON�iI M_IF1� D $ENA�BLE k LA�ST_^  d�U�K}MAX�� $LDEBU�G@  
GPCOUPLED1� $[PP_P�ROCES0 � �1��URE�Q1 � $�SOFT; T_I�D�TOTAL_�EQ� $,N�O/PS_SPI�_INDE��$�DX�SCREE�N_NAME {�SIGNj���&PK_F�I� 	$TH{KY�PANE7�  	$DUM�MY12� �3��4�GRG_S�TR1 � �$TIT�$I��1&�$�$T�$5&6&7&8&9'0''��%!'�%5'1?'1*I'1S'1]'2h"GSBN_CFG1 � 8 $CNV_JNT_* ��DATA_CM�NT�!$FLA�GSL*CHEC�K��AT_CE�LLSETUP � P� HOM�E_IO� %�:3MACROF2R�EPRO8�DRUeNCD�i2SMp5�H UTOBACK}U0 � �	�DEVIC#TI\h�$DFD��ST�0B 3$INTERVAL��DISP_UNI�T��0_DO�6E{RR�9FR_Fa��INGRES��!Y0Q_�3t4C�_WA�4�12HGX�_D�#	 d �$CARD_E�XIST�$FSSB_TYPi�� CHKBD_S�E�5AGN G�� $SLOT_�NUMZ�APRE�V��G �1_E�DIT1
 � Uh1G=H0S?@�f%$EPY�$OPc �0L�ETE_OKzBU�S�P_CRyA�$�4�FAZ0LACIwY1KR�@k �1�COMMENy@$DGV]QP� h���AL*OU�B? , $�1V$1AB0~ OL�U=R"2CAM_;1� x�f$A�TTR��@0AN�N�@�IMG_H�EIGHyAcWI7DTH�VTCYU��0F_ASPE�CyA$M@EX�P;$� Mf�C�FcD X $�GR� � S!1U`BfPNFLIC`~d
�UIREs3��AO}MqWITCH}cJX`N.0S_d�SG0� � 
$WARNM'@f��@� sLI? �aNST� �CORN��1FL{TR�eTRAT@0�T�`  $ACC�1"p '|�'r�ORIkP�C�kRT�q0_SF� �!CHuGI1 [ �Tz`u3IPpTYPVD�@*2 �P�`�� 1zB*HD�SJ�* ��q2�v3�v4��v5�v6�v7�v8��v9�vqO�$ <� so�o�h�s1��PO_MOR._ t 0Ev�NG�8`TBA � 5c���A�����]@B����ϋP�0XЅ*��h�`
P@�@�2� �,p�J,pC_Rrrqo@+�J/rL/�J�JVq@�Cj�`�m�g��ustP_}0sOF� 2  @� �RO_���WaIT<8C��NOM_�0�1�ەq3� ��cD !�;����hP���mCEXpG�0� F�<p%r
$TFx�J6F�D3ԐTO�3&@yU=0�� �YH�24�T1��E�� �e��f��f�>�0CPDBG;a� mk@$�PPU�3�f):��A��AX 1�dUN�$AI�3BUFuF��⠎�! |�`��`P�I��Pr�M�q�M~�䠁�Fr�SIMQS��G��Q�E������MC{�5 �$}1JB�`S��}1DEC�������ܴz� ě0CH�NS_EMP�r#$Gg�=Ǎ@_��q3�
p1_FP󔞡TCh�@`�b��q0�c}�y�G�� V�AԂ�!!���JR!0ԂSEGGFRA.pv 7aR��T_LIN�C��PCVF������Y ���Q��)B����( '���f�e �S���Q��.0�p�B�8�A����SIZC����z�T��g������QRSINF3��p�� ��?�������؉����Lot��G�*�CRC�eFCCC�`+���T� h��mh�SbA��h�*��f��:�D�d�c��C��PTA����w@��L����EV���jF��_��F��N&�G�� �X������1i��! ��,��h#RGNP��0qF���R�}�D���2}�LEW�N��Hc6���C�K�)�vqRcDx �:�L��ou2���A6N:`Co�$LGp���B�1aP��s@�dWaA?@���~0R���d�ME%`��d�_RAs3dAZC���z�OkqFC�RH`X`�F�`��}��,�ADI;� 6b� ��@�`�p�`5cn�S�@�1�7a�AMP���PY$8CU�MwpU��iQU� $�P��C��CG1������DBOPXWO����p$SK��2PP�]T TRL�1 ���Q0Ti� �P�DJ��4LAY_CAL`�1R !'PL	3&@�0ED�Q5'�Q5'"̡���1!�W�;PR� 
�1� 0�1" �PA�$�q$�� ��L�)#�/�#mp�0$��/�$C�!%�/�$E3NEqr�&�/�#�d REp�"'H� �O)@"$LF3#$�#xB� W;4���FO[ _D0m�RO(@���u��j��~�3RIGGER�6�PA%S���ETUsRN�2RcMR_���TU�`?�u0EW5M����GN�P���zBLA��E��$�$P#�CP� ��&�@�Qk�C5D�mpD��A#�p4\1i�FGO�_AWAY�2MO���fQg�DC�S_(<�QIS ����c�C���A����B�t�Cn�ȫA"�FW���DNT	V@��BVkQ�����S˳W�sU�J&�U�� ���SAFE�ZV_�SV6bEXCLUtl�����ONLA�b�SY��Q�tOTBa���HI_V/M�P�PLY_�a��VRFY_#�q�Bd��_ )0���_�+�Ip ���ASG3� *�b݀�0  AM���a*����0���Vi.b%fANNU�N� rLdIDp�U�2~S@�`mija�rj�f(�堫@I�"+���$FOb�׀O�T@w1 $DUMMY���d[!�d�١�& �E, ` 8�HExs���b�SB$�SUFFI�@ ��@��a5�g6�a!�DM�SW�E- 88�KgEYI����TMZ10^ӌq�1�vIN����q#�. D��oHOST? !�r ���t[ �t٠�tYp�p�EM>���$��SB�L��UL��/  �|3����T50�!?0 � $9��ESAMP�ԕF��׈�����I�0��$SUBe�Q�� �Cp�:��G�SAV�� r���G�C� ˇ�Pnf�P$80E��YN�_B�1 0�`D�Iad�@O���}�$]�R_I�� �ENC2_ST B� 2
ԇ J���L�@q~S�`;����!3��M�I��1:�p�4  L�3�M��0�0�K�4'a��AVE�R�q��}�M�DSP�v��PC�U��x�\ì�VALUŗ�HE� ��M�IP\@���OPP7  �CTHS ���6�S$�F�F􁳠dL�0�LT��SC�Q�d:��ETo�5zrFULL_DUY�da�0`��O�w�h�OT����0NOAUTO�!6�p$�\��R�cl�
�C` �IC���`!�L�� 7H *�AL���n�b���$�0 P�˴��ֲ��[!���a���Yq��dq��7��8J��9��0����1��U1��1��1Ⱥ1պU1�1�1��2
ʩ2����2��2��2�Ⱥ2պ2�2�2*��3
�3��3����U3��3Ⱥ3պ3�U3�3��4
�[�v��SE�"8 <��~��`�;I����׌/��QFE�0�0� 9� ,��Q? �z@^ ?�А��ER@#�`!�A��� �:�`$TP�$VARI�<��7UP2�P; �pq�TD��S|�1`3�纃�e�BAC�<# T�pr��)��b8P�P o�IFI)�P Ј������P�� ��0��� =t �;'�Ԡ��P'�ST (&�� HR&�r0E��*��	%�C��	��� _Cr�N�r��B��p�h�FORCEUP%b^n�FLUS�`H�N �E�h�RD_C�MK@E(����IN�_��&vPg�REMM�F~Q��M �� �3
K	N0�EcFF��N@IN�A��OVMl	OVA�l	TROV���DyT��mDTMX� ��m{@�
��? �*X[ ��CL��_:p�']@$�-	_
�;_QT��X
��@AQ	D� ��}��}!�V1� RQ��LI�MIT_�a椀�M���CLmd}�RIqV	�a��EAR��IO*PCC�����B�Bg�CM@��R{ �GCLF��G!DYM(/�aR#5TWDG��| s%��QFSS& �s> �P�a�!r1��wP_(�!�(�!1��E�3�!�3�+5�&�GRA����?w��kPW晅ONT��EBU�G)S&2*�P{@a�_?E @ �p�Q �TERMB5yAK5��ORI�G0BK5@�SM_ȣPr�G0CK5��T�A�9DK5� �UP>B�E� -zAa��@.PY3.@A$S�EG�:f ELEUU�SE�@NFI,���2�1ޠp4�4B$sUF6P�$��FQ4@�wAG0T�Q�&�HSNST P�ATm�piBPTH	J�AߠE�p��2�P@؀	E)�؁��1R�@<�InaSHFT_��1|oA�H_SHOR �ܣ�6 �0$�7�@Dq�'�OVR#�na�@�I�@�U�b �QAGYLO=�z��I'"��oAj�!�j�ERV ��:Qh��J��OG @�B�0����U>���R!P"�ASYM.�"��1#WJG�уES�A�YvR�U�T @���E)�ᥳEP!�WP!�W�OR @MB��GR�SMT�F�GR��3laPA.@��`|�q�uG � ����TOC�1�`P<�@ �$OP���P�pՓá ��O�񖌀RE�`RC�AOX�pтpBe�`RmE� u�h�A��e$PW�R�IM�ekRR_p�c4��qB H2�H���p_ADDR~��H_LENGqBPyqnq�q�R��S�I H� S���q0���u>Ӵu���u��SEȸ'�LrS��J� $N�`��_OF�F��rPRM� ���HTTPu_�H�K (��OBJ?"ip��$���LE`C!�ȠL� � �׬�AB%_~TS�s�S{`��6*�LVN�KR��e�HIT��BG��LO�qt�fN�͂���`���`SS{ ��HQW��A�M�p`�INCPU�"VISIO�����+��t�,��t,��� �IO�LN��N̠�C^��$SLQb��oPUT_�$�`�{�P �V���F_�AS�"O��$L ��I����A��U�0�@��af��`q�<PHY����Ó[���UO��#P `�����@�ڔ� �2�pP���`(�L��Y�B�Z�UeJ�Q�z�NEW�JOG-G��DIS�x�[�K-�f�#R �
�WAV�ǢCTR<�CǢFLAG�"[�;LG�dS ����Y�3LG_SIZ�o���������FD)�I�4�E�*�� D0���c$���𖶀����K���D0��� SCH_��߅p�2���N��F�T���E �"~�������U
�
�r{`L�	�DAU/ŃEA�-��dE�;�G�H�b9����BOO>��Uh Aɒ���IT��y�[0ŖREC��SCR��ʑ�DIēS.@��RG O���˒����d�´���SU���W�Ĳ��JGM$�MNC�H,�FNKEY�%�KM�PRGK�UqFY�PY�FWDYػHL��STPY�V`Y�@Y؀�Y�RS��H1`uۺ�CT���R��� �$�U	�m��� 
R�ݠғ`�G=��@CPOd�ڻŦ�M��FOCUd�RGE]X��TUIK�I{�����	������I�M��@A�S�`���@8������ANA���2��VAILl�CL�!�UDCS_HI+4`�s_�Oe�
!h��S���|�S����I�GN4��F�J��T��be�_BUj � Vj !PT�$*�@�rv�Ϥt���AVrW !Pi�'���0*�1?2?3?|_� X � i�`=a�5���Ņ�ID� tbP5R�bOh ��\AV�ST	�RF�YS0��@�  W$E�C�y����^�� Y L�؟0 ��@���`qFtǀ��FwҬ�_ Z i`����b���>0�C��[ �p CL�DP	��UTRQL�I{��T����FLAG�� 1�O�D������LD���ORG������hW>(�siT�r� 4\ ��#0��վ�Sy`T�70#0' �$�!�#RCLMC�$B/T/��)Q��!=1I�p_d]� d�RQ73$�DSTB�p�  � 6��-8AX�R |/8I<EXCES�b��2Mp�1^���2�Tt6��0_�p"6_A:&��;G?Y8�0K�d` \�G�ROU��t$MB� �LI9�CREQGUIRDB�aLO#KODEBUr� 1LYM��agbʑ`@�C�" 1ND��`c`ab���̨�CDC���IN'��C��Z`����H��N�"�a#�� �EPST�� cn\rLOC�RITp���P�Ap�1 �$��`AQ��d MX�ON�cF� R�fV�	X��b�U����uR�FX0IG}G�� e �y @X�a��X�XR�Q%��Y	��X	��V<�0ғDATA$`�E�a��a�N��f t $MDEaI:�)Sf��^d�![g�H5P�@]ez��a_cANSW�a^d�a��^eD�)DACPz�� nXpg �0CU4��V�`�=R0RR2�{�h D��`A��A��! d$CALII&0��GS�w2K��RINb�t<�NTEg�(i�bCu��X=RBqg�_N�qjPu�kr���$ht�2kuyDIV�&DHi0jp+�l $Vp�C�;$M�$Z0R<!�T 0R���b�em�H �$BELT|˪ZACCEL��q�;�"�IRCO��݁m��T���$SPSi0�Lt�ڰ�W��Cp8��T�9�P�ATH���.���3]��Pl1_<�r��Ł�"S Cr��_MG��$DD�9���$FW�`7`����.���DE�PP�ABNe�ROTS�PEEՂ@L� J�N�@��(0�t�$OUSE_p�P&�FܦSY>��p�! �Q�YN0A����OF�Fua��MOU߁N�GJ�܀OL~�ٔINC�d2Q��-2��<� -2ENCSpa`2U��+4R�IN��I]�B����"n�VE���s^�23_UP�օp�LOWL�� [�` '���D>�2 �PEp]'��2C[pW�gMOS���4MO���0�'PERCH  ��OV����蓼 ������$�8S+�� 2@������V�0^��O�L�P��7O�U�U�P"�������TRK|��AYLOA� J��1��]�͵³3P� ��RTI�1	�� MO�O�-2�28 �`4��wٳ��?�pD�UM2��S_BC?KLSH_C]�P� ϐΦ����bn�"�y�xÑ���CLAL �V��!��� ��CHKt �SՐRTY�� ��C�
*!6a_�ä'_UM����C����SCL�W�LMT�_J1_L< 0-օa:�E4�U�G�D�8J�P�J�SPCd�ȑ�Z���3�PC �3�H�_A@���C� cX�T���CN_rN����.�S��%�V ���:����]�9���C' �SH�r� *�*!9�9� p��^����9���PA���_P��_�"�Ŷ�!ճ����JG����~��OG��,�TORQU��ON��޹*�B0٢-�*�L�_Wž��_�sj��sj��sj�I*r�I��I�sFKP]�aJ�!��c!�VC�0'42��1��{0��82��JRK��+~� DBL_SM��:�"M�@_DL�q�"GRVq�j�sj�s�KH_��I���
CcOS��LN-  �����p�	�p�	�����FZ� ٦KcMY�D�TH��eTHET0��N�K23�s��s� C-B�CB�sC&1n2������s��SB8�s��GTS�1W�C.�2Q�����$�<'3$DU���8�A!r�2P&�1Q�b8V$NE�4�PI � ���"%�v$�p��A��%�'���LCPH�5�"h��"S�� 3�33�"+3:2�pV�(V�(�p�,UV�*V;V;V";UV0;V>;VL9H�(@�&�2�-n�H;H;UH";H0;H>;HL9�O�,O�(O}I�.O��*O;O;O";O*0;O>;O2F�"��Y�T�'SPBA?LANCE_T@S�LE�H_�SP�Hq�hR�hR3PFULClX�R{W�R3�Uz1i
�UTO_<����T1T2�Y�2N���`��Tq����Ps d���T�O��p!�L�INSEG���REVf��Q�gDIF��zy1j_g6�r1k��OBUa���t$yMI`���SL�CHWAR>��A�B��u$MEC�H�Tˑ�a��AX�˱Py��f�'�r�Pl� 
�bI��:�RO�B�CRW�-u����pMSK_KP�tn� P �P_��R ��r_tn���18�c��a�_p`�y�_p�aIN�:a�MTCOM�_C���po  �݀g`4�$NO�RES��r��`�r7p 8.�GRJ��e�SD� ABג$?XYZ_DA�!F�r�DEBU:a�q����pq _P$��COD�� 1����`���$BUFI�NDXa�Hp"�M{ORRsr $�q�U&���u��ӑy��^��bGi�s � $SIMUL���8��>���F�OBJ�EjP��ADJUS<ψAY_I��8��D���s�Ԑ_FIב=s�TZ��c� ���`b�"�(�b`p0:G�D��FRIW�d�MTg�RO%�A�Eb�z��HpOPWO> �Vpt0>�SYS�BU0[�$SOP���I�����U��b`PgRUN�rڕPArp�Dٖ�b��1�_OUbTΑ�a�t$�/IMAG��\pv �PDaIM��1�IN�[ �0�RGOVR!DY�˒���P�/�a�� L_�PB�}��¦�RB�� ��MLkᜪEDb��` �%N�@M��~���]��SLjPVpu x �$OVSLfS;DI��DEX���q �����o��Vb��N�A��'��,�'��D�M~��\�_SsETK�Vpv @.��^��ep�RI��j�
Bq�_�}����� Hp�dà*� w Hx\q�`��ATUS<�$TRCx T�X�NѳBTMڷıI���P�4}Ѱ���Vpx D\pE���β�0�Ehbϱ�����ϱEXEհ����)�=��bf�ym�]p԰UP��L�$�`6�XNN����������� �P�G�uzWUB�ñ�e��ñ��JMP�WAI[�P���L�O7��pFA`��$�RCVFAIL_Cwq�p��R9��p�c���(�}�"�-�AR_{PL��DBTB��,��pBWD ��pUM*�"�IG�7��Q�c�TNLW�"�}�Ry�iӻ�E�����Hp���DEFSP` �{ L\p�`��_8��Ճ��UNI�����Ѐ�RD��Rb _LA`Pͱ%�ѦpUq|-�#��q�O��XP:c�N�PKET�
���Pq�Uq} h~�ARSIZE5p���=��u�S̀OR~��FORMAT�P�g�COנq�<bEM2�d����UX��,�Γ�PLIb�Uq~ � $�pP_ScWI�`��IpAXG�~b�AL_ o�J��A�rB���C�r�D��$EL����C_lі� �� � ���r��J�30 �r��TIA4�Z�5Z�6�rMOM���f��s���pB��ADf��s����PU�NR����s������+��Rt�� A$PI�& E�kqE�p-~-� -�WC�0$��&��9q�gE��eSPEEDL@G���� �Ծ����)�9�����)��	)���SAM�WPx�0�1��MOVD�H$_S`Y%nk%$_��1�t�2�t�� ��c�v��8�H�PxIN����������(�+(+GA�MM<Vu!�$G#ETE�U�ٓD5�=
�PLIBRv���]I�$HIu�_L�HݰpB�&E�(A�.� �&LW�-�&�,�)�	6�&1��f�`j��� �$PDCK����ٓ_���� �E���b7��a4���a9�� $I
��R�`D�c�b~���`LE�qkq���81�¶0�����`Vp��P/aUR_SCR���A�r��S_SA�VE_D��8Ex�NO5�C��y�6�8@{$ E�.{I��G	{I�@�J �KP�q��H� ��� x"Mao���s� ���d��6W2U�Cq�y�Gq��M� � k�F��aE��3�W<�@[�jQWg@5r�U�RA�R��Sc2jQM"�&�[CL�W��M)ATr�� � $PY�����$W`�fNG�O�`�b�b �b#�HЈ��a� ���c��X�O���Zp�e��ހRt� p��p�3+zO�O�O�O��O�a5�_�r� | �E�8@��>vs�>v�� 8@_�kwVvy�Eހu%� C"rB�\�tP�"tP���PM&��QU5 � 8�*�QCOU�1 �Q�TH#pHOL<�Q7HYS��ESe�q�UE�p.BZ�O�䉋  q�P���%��U�Nְ�Q ��OE��p� P2�3��8AÔ�ROG����
�Q2(�O}�2�������INFO�q� �#�e����RȾ�O�I��� (�0SLEQ�с�рi�C��{�D��L��`� O�K0r��!E� N9U!��AUTTA�COPYqu�?���`@ML�NI�M�X�C�ᐛ� Y�RGAD�J�q�i�X�Q���$ഖ�`��W��P����0�������EX�8�YC0b�ѪO�bp�q���$�_NA9!�������`~��� � Q���POR�A�B��SRV0�)a�Y�DI��T_��{��������������5��6J��7��8y���S8BzL��m�MC_F�p
��PL9A8An�ȰR��9��Ѽ��$i�B����d� ,�0F1L-`L�C@YN�[��M��C?��PWR�c��L��!�DELiA��8Y5�AD�a���QSKIPN� �Q�4�OR`�NT�Q ��P_ 4��ַ@lbYp� ���������Ƞ���ՠ��������9��1�J2R� L��� 4*�EXs TQ %����(Q����p������p���RDCf�S �`��X9�R�p������r��A$RGoEAR_� IOT�2FLG��vi��M%sPC��B�UM_��~��J2TH2N'��� 1�����G:8 T00 ����ЉMlѺ`I�8��R�EFr1�q� l<�h��ENAB{�(cTPE�0�1��� i�m���^QB#��:��"P������2�ҙ��@��������&�3���7�I�[�m���&�4�қ�����������&�5�Ҝ1�C�U��g�y��� ��6�ҝ����������
&�7�Ҟ+=Oa(s�&�8�ҟ������&�SMS�K�q�|��a��E�?A��MOTEF����a@��(Q�IOQ5�Ic(P���R �W�0L�� ��pZ����#p%�L���U�"$DSB_S�IGN�1)Q%���C�l�(PeQRS232���b�iDEVI�CEUS�,R'RP�ARIT��D!OP�BIT`QY�OWCONTR;�(Q�ѬO'RCU� MDSU_XTASKT3N�p�[0�$TATU`P%�S�0L����p�_,PC9�$FREEFROMSp���%�GET�0�U�PD(�A�2%V"P|� J��� !)$USA^���6<���ERIO�P@&bpRY�5:"_>@ �qP}1�!�6WRKI�[D���6��aFR�IENDmQ�P$�UFw���0TOO�LFMY�t$L�ENGTH_VT�l�FIR�`-C�RSyEN ;IUFINR:]��RGI�1ӐOAITI��4GXӱlCI�FG2�7G1�0�Ѐ3�B�GPR� A��O_~ +0!�1R�EЀ�E3�e�TCp���Q�AV �G8��"J���u1~! � �J�8�%��%m��5�|0G4�X _0*)�L|�T�3H6��8P���%r4E3GU�W�P�W�R�TD����T���а��Q�Tm�$V 2����1��R�91�8�02�;2/k3�;3�:iva�9=i��aa�^S�jR$V��SBV�EV'�V�B
K�����&c�p���F�"{�@�2q�PS�E��$.rRC���o$AŠFwPR��Gv]U�cS'�� 7�8��E2I�� 0�@qV"`��p�d`���E0��@��=�
B5S!� ��aRg����iR�6�N AX�!�$�A�0L(A���rTHIC�1Y���h��t1TFEI��q�uIOF_CH�3�qI�G�a�pG1bxf����m���S@��_JFf��PR�ֱ�S��~Ԁ�d �$S�z��Z�GROU��̃TOT�t̃DSP�JOG���#��_P��"O������j��&KEP(�IR�����@M�R@�AP��Qn�E^�`�!�[�ScYS6��"[�PGu��BRK�B �.��pIq�p��M���΂�`�AD�!̃9�BSO�C׆�NӕDUM�MY14�p@SV��PDE_OP�#S�FSPD_OVR�=���C���OIR�CNm0�F.�l���OV��SFR��pU���Fn��!#��C8��A�"LCH����FРOV�s0��W�@1M��ĥ:�RO�#ߑr�_�p�� @@��u@VER�ps0OF�Su@CV? �2WD�6���2�ߑj2Y���T�R�!���E_F�DOY�MB_CM4�D�B�BL�b>�f��attV"Q�240/pd��N�Gg�z�AMx�`Z�0���¿_M~���"7����8$CA��7�D����HB�K81��IO�58���QPPA�=��"�M�5�͵���DVC_DBxC~� �3"�Т�!��1��糖�3����pН�*��qU�3��CAB���2VӆPѣIP��c�O���UX�SUBCPU�r	�S�P P� ��90^SQ׹c��."��?$HW_C�Т���S��cA�A�pl$�UNIT��l��A�TTRI"���	�C�YCL��NECA���J�FLTR_2_FI_�G(��9&�1�LP�?�>�_SCmT�CF_��F_�܌6��FS8!����CHA�1�wᇲ�"v�RSD�4"����qv�_T��PRO��,>�� EMy_ܠ��98d��a d��a���DIb0!�RAI�LAC��9RM��L!OÐ C��Q*q��X3q���PR��SQI�pU�Cr�s 	��FUNC��@rRI�N'PѸ0��u��!RA��B ����F��Ğ�WAR~���BLQ����A��������DA����	����LD)0��Q1�q��*q1TI2rQǁv�p$xPRIA1V�"AFB�P�!|�ߠ�<`�R���MO9I��A�DF_&@��l51��LM��FA�@�HRDY�4ORG�6 H���A�0 �MULSE&@"�Q��a� �G�	������$d$�1�$1 ���0���o� xm�EG�̃�`ARހ���09�2o��z�AX]E�ROB�W�A2��_�œSY���t���S�WRI�@rs1��STR��� ��(�E�� 	%1��AB( �/&X�a�ӰOT0^�;	$ߠARY�sf"h���S@	�FI��~*�$LINK����!�a_%#�t%{q�"XYZ828�*�q�#OFF���")�"�(j B�j��4С��n�3FI���%7�q���j���_�J���%��#�QOP�_>$H+5�3�PTB�\1�2C��i�DU��&62�TURN ��2r�5t!}��p��|7FL�`���m�0�%�+*7�	� 1�J. K�M�&82�pQ�2rQ�#�ORQ�� G��-(�+p��z�� �3q�E"��T�GOV�@-A��M*�y�4�E:�E@�FW�J��G ���D��o�*� ��A 7�P��y��E�A�GZU0:ZU�CG�ER���	6�E���B�TA FQ��)4����r'�AXУa2.q�c �W�c�W�c�W�p�Z�0 �Z�0�Z%@�ZK@�Z� �Z
!�V� �Y� 
i�  i� *i� :i� Ji� �Zi� ji� zi�a�iD7EBU{�$v�u���;q��"F7O�n�A!B��6��CV�z� 
fr����uk� �w�!�w�!�w�1�w�1 �w%A�wKA�w��\0���"3LAB"2�|EwЄ�҂�3 } EERVEN�� � $q�_NmAǁ!_�PO�����` f�M�_MR}A��� d  9T���ERR�����~ TYi��RI�V8"0�S��TOQ�T)P!L��T�ЅL�G�}CJ � p�PqTl X���_V1�bP�Q���#�2�2+������/@��p��5��$W��V���VN�[�$�@�� �S����Q�	EHELL�_CFGN�� 5%�B_BASƴ�SRvp0�K� E�S��Jϐ1a�U%Α2�3�4�U5�6�7�8�RO���� � NL:�3ABn��АACKwv��)�o�pu0iႩ_PU2��COq��OU��P���ӕ�����T=P�_KAR�0&��REm�� P����QUE٩��@����CSTOPI_ALzs��� �T���� SEM[�w�k��Mw�y�TY��SO`��DI���Є�=��װ_TMK�MA'NRQζ� E���$KEYSWI�TCH��Ѱ��H=E��BEAT���EpLE����&�U���Fd�����SO_�HOM� O��REF�@PRi��R� ʞ�C@�O0�p EC�O���� _IOC1M�4M�k�L���'�O� D�!ۧH�	U��;�M7��@�3�FORCߣ�� �_��OMq �� @Etxk�U#P�o1B�O�o3B�4�x�NPX_AS� 0ݐADD|��(�$SIZߡ�$VAR�TKIPr�q�G�A(����
�˨r�t�n��SV�XC����FRIF�R��S%�7�xĆ��NFѲEАO�� x�PSIڂTE�C*�%CSGL=�T�"�0&�V�D��>�OSTMT
�o�P\��BW�@?�SHO9Ww��P�SV� K߹� ���A00�0�Q��K���O���P_���i���5��6��U7��8��9��A�� ���6������20��F��
 ����U ���� � ����0�� �J@���:�1G�1T�1a�1�n�1{�1��2��2���2��2��2��2��2�2 �2-�2�:�2G�2T�2a�2�n�2{�2��3��3���3��3��3��3��3�3 �3-�3�:�3G�3T�3a�3�n�3{�3��454���4��4��4��4��4�4 �4-�4�:�4G�4T�4a�4�n�4{�4��555���5��5��5��5��5�5 �5-�5�:�5G�5T�5a�5�n�5{�5��656���6��6��6��6��6�6 �6-�6�:�6G�6T�6a�6�n�6{�6��757���7��7��7��7��7�7 �7-�7�:�7G�7T�7a�7�n�7{�7���+���P$�UPD��  �P���x��YSLO��� � ��հ�����Q�TAS�sTƠ��AL1U}U����CU��W=FdQID_Lѳ�U�HI�ZI�$FI�LE_Σ�T�$�u�_VSA��� h���+`E_BLCK�(�8bg�AhD_CPUQi��Qi���Sodx_R1�ɢR ��g
PW,�d� �aLA�S���c�a�dRUN5��a�d�a�d���5��a�d�a�d ��T�pACC����X -$&qLE�N~�3t��&p����I�ѱ
�LOW_AXMI(�F1&q�T2mwAM��ɢ����I��8��Q�yTOR.�&p�{DW��s�LAC�E���&p�����_�MAuйv�u�w�qT#CV�|��wTڱ� ;�1�<ѷt��_��s��IJ����M��ӠJ�����u���u2q2���������s�pJK�цVK~�か��3fՃJ0���JJ�;JJ��AAL��(���4�5Xr;��N1B�N��	��tL��p_k��?Q"p���� `5`GROU�PY�ӲB$�NFL�IC�ө�REQUwIREv�EBUV�0"q���кp2���#p�ɖ!qxг�� \^��APPRՐC��ڜp
!�EN�CL9Oz�,�S_M ����A��u
!q��� 䣠MC�r;�Xr|�'_MGц�C��,`p��N��p��BRK��GNOL������Rϰ�_LI��է����JޠѤP��p��p�� �p;��pD��p6�K���8��n�"q���G� ҒMr:ql�<Gqz�PATHv���@����Rx�������pCNR�CA��է�6��IN%rUC�pwQZ�Cd�UM�Yop�����QE:p�Gp������PAYLOA�ͧJ2LHPR_A	NqQ�L�`[�W�K��g���R_F2LS3HRё�LO\�������ACRL�_�����޷C�XrH��P"�$H���FWLEX� qJ%u� :2Dv�p 4�K�GYq�pPbt|F1Kљխ׃�������E��� �/�A�S�e�w����� y���ф���蘏����$J�ÊT���X���� υ ��څ��[���� 
�� �)��;�D�V��h�z���J��� �� �������QIPA�T��ё��EL4� ��ؘJ���ߐJ�E��CTRޱ��T�N��F�ɗHAN/D_VBp�ѹPn`�� $&�F2��XK��ШRSW��Y��j��� $$M��}�R��E��Uw�H��sA�PH����QD���A���P��A��AAɫ���j`��D���DɫP��G�`1)S�T��9!��9!N̨DY�`���|�Y�� ��KыǦ�J�ч�s�U�ХP��&�/�8��A�J�S��`�� �; �t�.R66N�/QA'SYM����Ґ�����Խ��ٿ_SH �����筈4��+�=�O�JV��h�'C�I����_VI��dHN�u@V_UNI�ÉD���J҅�B�% �B�̦D�ųD�F�̓�@�������*Uc���ӆ��H�`���XQEN� v�DIɠS�OwTY�YP���� ��I�1A ��äQ�`Bc�S`� � p�a.a� � ME����R'R�1TkPPT�0) ���Qz�~���0�Xa�	iT@� $�DUMMY1��o$PS_��RF���X�$Pf�aLAƏ�YP�jb�S$GLB_T>mU�e��PpQ p���Q� �X	�ɗ`�ST���ߐSBR��M21�_V��8$SV_�ER��OÐ�c�cC)L�`�bA5�O�RTP�T O�P � D� �`OB���LO˰&uq9c�`r�0�SYSqADR��TP�PTCHb �� ,&����W7_NA���tz�삑Y�SR���l =��M�u` �ys�u~�s��s� ����������0� )�T�"�5�~���B�����s�?�?�?DY�XOSCRE)�p��ȐST[�s}H�P!��t�Qr _� Aq� T	��`ob ��a`�l��Ҥ��g��c�O� IS��c��UY�UE�T� ��ñjp^`Sq�R�SM_iqmUUNE�XCEPlV֑XPS_�a����޳����޳R�COU�ҒS�o 1�d�UE�t�ҘR�b9�PROG�M� FL�$C�U�`PO?Q�д�I�_�PH�� � �8џ�_HEP������PRY ?���`Ab_�?dGb��O�US�� � @��`v$BUTT��RV`��COLU�M��U3�SERV<x��PANE� qu��P@GEU��<�F���q)$HE�LPB�l2ETER��)_��m�Am��� l���l�0l�0l�0�Q�INf��S@N(0�� ǧ1����ޠo �)�LNkr'� ��`T�_B����$H�b TEX�*��ja>�REL�V��DIP>�P�"�M�M3�?,i�0ð�N�jae���USR�VIEWq� <Ե`�PU�PNFyI� ��FOCUPn��PRIa0m@`�(Q��TRIPzq�m�UNP�T� �f0��mUWARN|lU��SRTOL�u����3�O�3O;RN3�RAU�6�9TK�vw�VI͑�U�� $V�P�ATH��V�CAC�H�LOG�נ�LIM�B���xv���HOST�r!��R��R<�OBOT��s��IM�� gdS X`} 2����a���a���VCPU_AVA�ILeb��EX��!W1N��=�>f1?e1L?e1 n�S���P�$BACKLA�S��u�n���p� � fPC�3�@$�TOOL�t$n�_wJMPd� ݽ��U$SS�C6�Q�VSHIF ��SރP`V��tĐG�R�+�P�OSUR�W�PRADI��P�_cb���|a�Qzr�|�LU�A$OUTPUT_BMc�J�IM���2��=@zr��TIL��SCOL��C����ҭ�� �����������o�Bod5�?��Ȧ2Ƣ��0�T���vyDJ�U2��� �WAIETU����n���%��{NE>u�YBO�� �� $�UPvtfaSB�	TPE/�NEC���  �ؐ�`0�R6�( �Q��� ش�SBL�TM[��q��9p����.p�OP��MAS�f�_DO�rdATZpD�J����Zp��DELAYng�JOذ��q�3�����v0��vx��,d9pY_ ���	�7"\��цrP�? O�ZA;BC�u� ��c"��ӛ�
  �$�$C��������!X`�P� � VI�RT���/� ABS�f�u�1 �%�� < �!�/�/??0? B?T?f?x?�?�?�?�? �?�?�?OO,O>OPO bOtO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_�_�_�_�_�_ o o$o6oHoZolo~o�o �o�o�o�o�o�o{� >��AXLMT�s���#  �tIqN&8qtPREO���+vupXuLAR�MRECOV ��)XrzujF }�%�!d�������7�I�[�m�~�, �
�/��vNG5� ��+	 A  � ڏ�� PPLIMC5�?�%upՁ�Handl�ingTool �-� 
V7.7�0P/36뀬��
]�_SW2�D�Fy0j�W� 43Y��J�9�K�7DA7�?����
&�X�e�	-�None���J����� �T7��	���_�V�iu�6s��UTO�z"�,tTy.�HGA�PON� %��!.�U���D 1�y� t�x�����y.�K�oQ 1�{  Hp*������	����uq��"�" g�!��Hե�w��HTTHKY��"ٯ����u� ����󿽿Ͽ���� �)�;�M�_�qσϕ� �Ϲ���������%� 7�I�[�m�ߑ��ߵ� ���������!�3�E� W�i�{��������� ������/�A�S�e� w��������������� +=Oas� ������ '9K]o��� �����/#/5/ G/Y/k/}/�/�/�/�/ �/�/�/??1?C?U? g?y?�?�?�?�?�?�? �?	OO-O?OQOcOuO �O�O�O�O�O�O����TOĀ��DO_CLEAND���{S_NM  ɋ����_�_�_�_o��_D?SPDRYR�_��HI!��]@�_}o�o �o�o�o�o�o�op1CU��MAX � bTQNQS�sqXbTB��o�B���PLUGGpb�cWo��PRC4`B�P]klo^�r�O�r=o��SEGF;�K�+�6��_�_}��������ŏ�0�LAPZom�/��+�=�O� a�s���������͟ߟ|�6�TOTAL�v|�y6�USENUZ��g� HXL�NR��R�G_STRING� 13�
�kM,�S�
���_ITEM1��  n󝬯��Я��� ��*�<�N�`�r����������̿޿���I/O SIG�NAL��Tr�yout Mod�e��InpB�S�imulatedޕ�OutT��OVERRW` =� 100��In� cyclHŕ��Prog Abo�r^Õ�>�Sta�tus��	Hea�rtbeat��MH Faul����Aler���� �'�9�K�]�o߁ߓ��� ^S��^Q�� ������,�>�P�b� t��������������(�:���WOR 9���r���L������� ������*<N `r�������PO������ �9K]o��� �����/#/5/�G/Y/k/}/�/DEV� -�/�/�/? ?)?;?M?_?q?�?�? �?�?�?�?�?OO%O>7OPALT��^A ��8O�O�O�O�O�O�O �O__(_:_L_^_p_��_�_�_�_�_LOGRIxp��avO�_*o<o No`oro�o�o�o�o�o �o�o&8J\n�_*�R�ݦqo� �����(�:�L� ^�p���������ʏ܏�� ���PREG bNK��$�r������� ��̟ޟ���&�8� J�\�n���������Ϳ�$ARG_r�D ?	�������  �	$�	[��]���.��S�BN_CONFIOG ��L�K��F�CII_SA_VE  �k��b��TCELLSETUP ���%  OME_I�O��%MOV�_H��¿ȿREP��|��UTOBA�CK��V��FRA:\8�c �8���'`��q8�c�,�INIa@�8�^�,�MESSAGz������>��ODE_D��}��C���O� ��,�PA�US!��� ((O��J�\�F� |�jߠߎ��߲����� ����B�0�f�t�%�~*TSK  5�x�ϕ�/�UPDT����d����XSCRDCFG 1��;� �������&�8�J�\�n��� \�n���������� "��F��j|�����/e�2�GR�OUN����UP�_NAܰ��	�2��_ED��1
���
 �%-B?CKEDT-���}��pg���Pg3�p8�/�/�8���g2���E/��/��/~/��ED3n/&/�/J/�\.�/"?�/�/ED4 ?�/?�/\.[?�?5?G?ED5�?n?#O�?�\.�?jO�?�?ED6 ZOO�O6O\.�O_}O�OED7�O�Ok_�O�\.G_�_!_3_ED8�_�o�]-�_Vo�_�_ED9Fo�_�o�"o]-�o�oio{oCRoY_Vh�]1��{� LNO_D�ELGE_U�NUSE	LA�L_OUT �V��WD_AB�OR���~�5�IT_R_RTN�ǀH�ONONS)Ю������CAM_PAR�AM 1����
� 8
SONY� XC-56 2�34567890�Y �f�@����?�W�( С���8�h�х�ڎ��HR5ǃ��	���R570�B�Affފ������ڟ� ǟ�"���F�X�3�|����i���į!�CE__RIA_I����5��F��;�Я� ���GP 1]����s�����V�C󠸾�����CO�C ��(���ǀC8��@��H̺�CCX����Ch꺰p��x���� +C�����Ⱥ���+�=�G��ށ��HE>/pONFIG=�f��G_PRI 1�B�$r�����������(�~�CHKoPAUS�� 1���� ,wuj�|ߎ� �߲����������� 0�B�T�f�x����D�O���T���_MORGRP �2?� �\�� 	 �,��P�>� t�b���5�����eҒ.�?a�a�����K(���d�P�V��a�-`�/A�

s��������b&�i��ܦP�DB�����)
�mc:cpmid�bg��:� � �+����p��U   ��  �s�3�� ��dܷ·{C�e�*����{g�+/*���{f/s/�i�u/�
DEF ��(K�)�b b?uf.txt�/\�/��_MC����E�d,53������ʇ�Cz  B��p�B�Z�B���B�;@B����B��
C3�"
q�Dv���D/DF���DRt�DC$�D�QГ=F�p�gF��FM�F�EF�2�?FLE�	?B���
5����S4���(D~���/�v̂3@�à1/  TB�D=�V@a  EI�5�� F*� F��G$ˀF[�� GR�kNGl���G��G���&H��G֓ϦH��߃]�� � >�33 9�ށ�  n^���@߂5Y�Ed��A���=L��<#�
 ��_�*~2RSMOFS���.^�9T1��D�E ��l 
� Q�;�P  x0_*_>TEST�")__��R���#o�^6C@A�KY���Qo2I��BR ��� �C�qeT�pFPROG %�(S�o�gI�qRu�����dKEY_TBL�  6��y� �	�
�� !�"#$%&'()�*+,-./01���:;<=>?@�ABC� GHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~�����������������������������������������������������������������������������q��͓���������������������������������耇���������������������9�Eъ`LCK�l��<�`�`STAT�c�_AUTO_DO���O�INDTO_ENB;���R�Q�Y�K�T2����STqO�~��TRL�`�LETE�ފ_�SCREEN �jkcsc� 	�UπMME�NU 1i  <�l�ol� K�u���FS����柽� ϟ���R�)�;�a� ��q���Я�����ݯ ��N�%�7���[�m� ������ɿ�ٿ�8� �!�n�E�W�}϶ύ� ��������"����1� j�A�Sߠ�w߉��߭� ��������T�+�=� ��a�s������� ����>��'�M���]� o��������������:#p)+�_M�ANUALӏ��DwBCOu�RIG��$�DBNUMLI�M�,1e
�P�XWORK 1k�_-<_N`�r�TB_� � m��Y0�_AWWAY��QG�@rb=�P�_AL� =���YҀ��`��_�  1!�[ , 

:&d2/(o/�&�Mt�IZP��@P�#ONTIM6��d��&��
�e#MOTNE�ND�o$RECO_RD 1'kU2)?�!�O�?1-?&k �k?}?�?�?88�?�? ??�?c?O*O<O�?�? rO�?�OO�O�O�O�O �O_�O8_�O\_n_�_ �__�_%_�_I_�_o "o4o�_Xo�_|o�_�o �o�o�oEo�oio�o BTfx�o�� /�����>�)� 7�t�� pu�����-� �͏ۏ�����N�`� Ϗ��o����)�;�� ����8���\�˟ݟ ����;�Q�گI���m���4�F�X��TO�LERENC�B��	"�L�Ͱ C�S_CFG (� +x'dMC:�\��L%04d.'CSVY� cֿx#[A ��CH�z _/x.�G��},���RC_OUT �)�- z/��SG�N *��"���#�27-M�AY-25 18�:41����4:�38�]� Z�t�����x.�����pa�m��P�JP��k�VERSION ���V2.0.1�1~+EFLOGI�C 1+� 	d��ٓ��p��PROG_ENB��2��ULS�' ��p�_WRST�JN� ��"�EM�O_OPT_SL� ?	�]�
 ?	R575x#?�74D�6E�7E�50i�d�o�2E�d��|j�"�TO  .�����k�V_� EX�d�% �PAT�H A��A\p��M�_�~+ICT�-F�, '�`ßeg��}�STBF_TTS�(@�	��Eм`���� �MAU��ߧ"MS%W��- )��},t�
��.�!��]l�R �v�����4�SBL_FAUL�y�/��#GPM�SK�ߧ"TDIAb��0����`���!�123456�7890xS�l�P �����//%/ 7/I/[/m//�/�/�/��/�/L0PV ���/�2? X?j?|?�?�?�?�?�? �?�?OO0OBOTOfO�8<x�UMP$�I� �ATR>�Oδ@PME���OY_�TEMP��È��3��4��DUNI�	�w�YN_BRK� 1��x�EMG?DI_STA	���GUNC2_SCR 27[��_�_ �_�_�&�_�_o o2or�nSUQ13y_+?|o@�o�o�olRTd47[�Q��o�o���_ >Pbt���� �����(�:�L� ^�p������� ?Ǐُ �0�,p��+�=�O� a�s���������͟ߟ ���'�9�K�]�o� ��������ɯ���� �#�5�G�Y�k�}��� ����ſ׿����� 1�C�U�g�yϋϝ�ׯ ��������	��-�?� Q�c�u߇ߙ߽߫��� ������)�;�M�_� q��ϧ�������� ��%�7�I�[�m�� �������������� !3EW��{�� �����/ ASew���� ���//+/=/w a/s/�/�/�/�/�/�/ �/??'?9?K?]?o? �?�?�?�?�?�?�?�? OK/5OGOYOkO}O�O �O�O�O�O�O�O__ 1_C_U_g_y_�_�_�_��gETMODE �15'Efa �t|�_GgRR�OR_PROG %�Z%���Hog�TABLE  ��[1O�o�o�o�ZR�RSEV_NUM� �R  ���Q�`a_AUT�O_ENB  �u�SZd_NO�a �6�[�Q�b W *�6p�6p�6p	�6p�`+5pOastHIS�cXa�P{_ALM 17�[� ���6|6`+t���&�8�J�rx_�bp  �[�4q�R���PTCP_VER !�Z�!6oZ�$EXTL�OG_REQ�v9�y�SIZ�܄�TOL  XaD�z�r�A ܄_BWDo�%��fQ���w_DI?� 8'E�t�TXa b[�S�TEPg�y��P��O/P_DO�v$v`�FEATURE �9'EQ��Q�Handlin�gTool � �DER En�glish Di�ctionary��7 (RA�A Vis"� M�aster����
TE0�nalo�g I/O��p�1
0�uto �Software Updateb�� "/�k�mati�c Backup~
�d
!���ground E�ditB�  25�LCame�raT�FX� "L�o��ellT��Lw, P��omm9��shۡ�h600���cou���uct���p�pane� �DIF���tyl�e selectvѡ- /�Con��~9�onitor���Hd�tr�Re�liabT�ϣ(R�-Diagn�os��Q�	�H�Du�al Check� Safety �UIFc�Enha�nced Rob� Serv��q ��v	ԸUse�r Fr���T_�i�xt. DI[O f�fi�� )��\�endܰEr�ru�L��  pr$נ*�rO�� @����ENFCTN_ Menuİv��.fd`�TP �In?�faco� � 
E�G��p;�k/ Excذg�C���High-Sp�eܰSki��  �Par+�H���m�munic��on�s��\ap��ur�f�?�X�t\h8yU���connZ��2Т !�Incr��str)�8���M-6�KARE�L Cmd. L���ua��}��B�R�un-Ti�En�v�(<�@�I�<�+���s��S/W�"�H�Licen3se���� ad����ogBook(S�y>�m)	���"�MACROs,~��/Offse\��f����H�!�Y�M�1�MechStop ProtZ��3� 5
�Mi�4�Shif\��B;6S�MixܰQ�����H�Mode �SwitchY�M�ok���.�� ��MTt�Q�g�� �5��?ulti-T����ܖ�)�Posj�Re�gi>���  ! ��PA�t Fun<1��6iB/��R��Num�Y�3�G�P�/��� Adju<��	�/2HS�)�� o(�8�tatu����AD ��RD�Mޱot�scove&� #e�v������uest 867.��o�\���?SNPX b��Y�<��)�Libr%�
�Ort I���� "����.S�o� ��s� in VCCM,����� j������㣀/I�� 7�10�TMILI�BX����g�Ac�c����C/2�T�PTX�� �Tel�n��Y@����K�P�CUnexc�eptܰmotn¾� ������\m725����w�|5���  h640SP CSXC��i � j*�� RI�N��We���50�,��vrl�زmcen" ��fiP-��a���P��Gri�d{�play F� O/��? ��EL�R;�|�20��O{RDK�sciiw�oload�41d�;st�Patd���CycT�h���or�iɰ:�7c DatMa� qu6�2�0��*�������FRL�amc�K�HMI De��(����k��PC�φ�Pass�word�644���Sp�����D#Y�ELLOW BO��	?1�Arc%�v�isu����#ti�O�p�^�! 2��a6O�po�� t��ֶcT1o�����HT���xy�	�  5 $�t۠ig��1�0Ơ 41\+�J�PN ARCPSOU PR+�8b!�OL0Sup�2fil� �!��E@-�;�7croc�82��v����$ 12jSS�0e4�tex-� �I�7�So��tf�ssag�� e��У�qP��,��� "Tc �Virt��v�!�����dpn�
�J�3�SHADf0M�OVE T�MO�S O TԠ�get_var ?fails l�>P�U~1E���� Hold Bus %��h��VIS UP�DATE IRTORCHMA A�|{�vYWELDTV �S ]�DtS: R�741��ouiPb�}�y��BACKG�ROUND ED�IT "RC$REP�TCD CAN �CRASH FR�VR 62z1�SC�ra��s 2-D���r ) "��$�FNO NOT {RE��RED �`� m ��JO� �QUICKaPOP� FLEN m4�1S�Loc��gRT�IMQ%�#�FPL�N: FG��pl �m�r`�MD DE�VICE ASS�ERT WIT gPCV;PB�AN#a�ACCESS Mo .pc��Jo���Qui±�Kbld�mgUSB$ ��t� & remov� Pg�SMB �NUL� ;a|�FI�X��C��ACHI�N,QOL�`MO �OPT ՠa��P�POST0�WDUs C�wQAdd�`�ad���0io�2֫�$P�`W\0.$�0`O�IN&�P:�fix CPMO�-046 isskueC�J/aO-�0n�r130Т- ���vRSET VAR?IABLES-P{�ޯR3D m��vi/ew d��M��&��ea���b��of� FD�5P:N@x� OS-1y0`�h� sc���t��s ft�lo��7 WA�P�Z�3 CNT0 1T�/"�ImR�)��ca �Pu��PO�T:Whenape=wB�STY E�{1�t��ptKQdo /GET_�p �p��VMGR LOl�REAd0C~QW�~1��(�l�s�gD�EC�TpLpING /IMPR�DR(p+P�B�PROGRAM��ERIPE:ST�ARTU� AIN�-;�ӠM/ASC�IIzPÂOF L�q�DPTTB: �N�pML$me hP���`:x�mo&��allW`!�ӤTo�rc�A�U�HC�i�LpԸth�`n�@ �ch��/GEA�!�t�ou͐�RCal���k�Sign`� �ND�ԗThresh123��`��09p� : MSG_P�+0er  �Q�=Aܠzeron���0 H85��RI�mA�n�2D��rc:�0I��OMEa`�p�ONaP5�  נS�REG:FF-Д� �]�'���KANJI*��n��J��c�0as�n d�!OA im�mc �INISI�TALIZATI����~1wem�����dr+� LB A|�UWqminim�rec[�c!�R���}m$�ro -1>��S�ܰir��@ұJ�*1pdETw�� 5`?��I�ow u��< s_e 1lc��YbPM���p�Q���R`vR�&�lu\�3�Re �0�4q�q1#���m9 <a�arn���~��Box fo���*PRWRI�PW�S���v�09 F�pu�p�de-rel2 d�p� j��`━�betwe��IN�D Q���igE osnap|�us��spo TME��7TPD#�DO�p#a�HANDL 1\�k�`vR��ȀD�n�y�S�v�Yoper�abil� �T*�:� H � l\p��V�q�b�R�< p�a*�c&2O�`FA,�.�-QV7. f.v��[GT�pi�s���� ɠtmLin�e-Remark� �� RM-�` �W�#SPATH S�A+PLOOS U�IFc�+5f fig��pGLA����Vrp�������U�0the�r�V� TracD���tW�\b�s7���d�t�� n�@ I ���3:���dK�=y��it k8�d�wPayR![2]��^�1: g��s���dow�XQ��0I�S�q�qEMCHK EXCE C����MF +�Xah>�� 35\k��)���QBt���'b�d��[�c���e �`xk�S�� BUGrt��cD$`PETpȵ��f�c4��0XP�ANSI��DIG���@OoPmetTC�CRG EN��C�EMENT�A M�̀K {�`H G?UNCHG �`� �EXT�P�2�bQS��93 wP8�x�O�RYLEAKq � H5gyq�PLC WRDN R �sO /u�QSPE=p��G*�V ��$��tn720\3pGR�I��A�rT�PM�C ETH��pSyU7p�`  j5/^n�PENS�PN,���*P ont�`B�ROW�`!sRMVo ADDz CN �qDC���PT3 �ALA2@ ���pS�VGN EARLqY�R��ŰH57�GaJLAYҀEk (@M�PPD�p:*@H�S I`P��OUCH8���V�F�q�comH�x ���ERROR� DE� nJ��RO�C�URS8pI��Nx4q�-158n7��RSR xP#aU�p���Rqy�T�F�z�;�pk��t�� �gՂ�B�SY �RUNN�  a|�`�BRKCT�!�RO�p3@ \ap�SТ�AXxP���h�8+ q��ISSU�r} sPX�PTSI��K1M10_�I�PSAFETY Ck�ECK[��Á ������<#X�� ��TWD2�@�@�I{NV��D ZOp�5X��t�DUA=Ly� "M6�0�J"rF#�E��dPd?NDEX F�,t*UF�"Pʀ��0sFRVO117� A�PT6�KtqF�ALPTP247�7D6_�P�!;HI�G� CC�t;SNPX� MM��tq�d~�Vq�q#�
"��>DETEC�Tq*@RRU�qA�P�5p�9 y�)<9���7T��Pds� k�	���!Q���� t\4A�;A0�o2 "Ke@" 8@�HI�qXF8@4@H�PRDC"�
�aMB8@�IXF�b���zOX@8@����a�G}E�B�Ccs�cr�J8@�Ndctrld.�A�NZE�A�5��Q��!�`�Df�8@�`m�878�Q-z;� ��� rm`�i
��PR̠78�@�RI8@0q�Q ( ~\Mp��0t��!{B8@�\tQ<OX�St0�32hB3nO�Vtp�A�@gLCF�L��� �Rplcf���J8@�WTamai�E8@mubov2_miTA�O�S8@�U`T[tT�AqPr67�4xSShape GGen��8@j�I�[R�`�@8@T����%qc (u8@��II�^��Q~C�a�[8@;Ynrsug0�4� � 4�C�tMr68@�r5hB5��zVnretsp e"r�Po�wng0bGCRE�Ka�ޠ��DAT�E�k�creat.�q�M��a�oksqgtpa�d1P��(�tput�Zj�{�������܆2�8@����Q����sl�o��� �hex�H�TB�8�ď�ke1yH�8@�pmZb�NbR�u7A+�nrgc8@ UQ�pp�bUZ�dp0a�j921xSpl.Collأcq�\A�b�RNq�UA� (J�8@ip�_�WA��_�Y���a7hB7�ͦt�p[� "TCLSx9oKb��clskyht[��s�pkckZd ���$�TQ���dA�r�x�710a- KA�REL Use {Sp�FCTN9��a�7l�0s0a�� ( ���a��~C8@��MI���c8hB8"   ��8@ v	��v	   �lmatea99�qM����E�mcc;lm5�CLM;�� ��j��E�et���aL1M	�h�yasp,���?mc_mot�B�N���8@H����Q��su�'��Q�ȕ�䅮���j�oi#�ߕ��A_l�og�Z���trc�B����ve�ϓ�v���QWX��6�find�erxSCente�r F1�lSw52a0��ha6rX� (<�cr,�Q�Ձfi�Q  �NH0�I�ۡ���A8@�uL��tq�a "F�NDRVϳ���et�guid�UID �C8@���������TA@�nuf;��P�����C�B��_z�Ӡo��qG������l���f�ndrTY��2䁴t�cp"�,qCP MtF�}38@517��6s38�E��gf6 ��(��K��Q��-�X�L�A�tm6�P�� ���Q���	�����tm�Ĵ�b8@aej��TAiex���aP�Aa�ذ�cpr�m�A��l�_vars��
��dwc7 `TS��/�6��ma7A�F�Group| s�k Exchan�gJ 8@�VMASK� H5�0H593� H0aH5@� 6V� 58�!9�!8\J�!4�!2���"(�/���;OMI� `@a0�hB0�ՁU4U1#SAK(x2�Q�0I�h�ӂ)�mq�bWzR�D�isplayIm�Q@vJ40�Q8aJ�!(P��;� 0a���0��� 40;�q�vl "DQVL�D쌞�qvBXa`�uG�Hq�OsC��avrdqq�O�xEsim�K�40sJst]��uDd X@TRgOyB�Bv40)��wA~���E�Easy� Normal Util(in��K�11 J553m�0b2v�Q(lV40xU�)��������k986#8Uϕ�|�rP "NOR��dw d.a}oKksu�O�W����OY�W`�j0�6�H� �menuuyP6�Mx�`wRX�R577V��90 �RJ989F}�49b\�`(�fity�����e��<?��Vsmh`��8@��C0�Sv�q�8����w�pn "MHMN<��ޣx�Ay`�o��3�u�`f�І�x�t ��tRzQ��LV��vP�#tm���|I�1{oPx" �2|���I�3I/B��odstǏًmnx����}ensu_�	L<���h!!��Rt~��huserp��0Ҹ�ʐcM�_l�xP�oe��рpoper�����xdetbo /�l>�x���Ps$p��`���OPydspw�eb͓��z'R��u�Rr101&S՟{tb�`2�Z4�30������`4�
�4�5���KQ�m[T��dUCalG40`�Q)p40}������9;��DA��? v	LATA�umpd�\bbk7968��68c�f�bl�41969y�9и|�D���bd� "�BBOXêM��s�ched����m�s�etuM:�����ff���40��n�41��8��40q�col��|��1�xc�ؘ���li ��X�0���j��&�8��4 <�ro5�TP �E�#��ryK412r��;�(T+Q �Rec'�ʈ1Iw��84�����Ak97�1��71�;���p?arecjo��Q�NS�[T���dXra{il| nagek��M ,QT2 *� !(�ĜR%<x�80P!bh��p��4���4�yDgl�paxrmr "XRM�g�l�brf{���n���kl��9turb�sp��㧑- �l0s15	�g�625C� Mh�+���)89��	+��B6��o�ҹ��x�7�q40�����pd "TSPDx�=��tsgl��l�:dQ���8Bc1t���K�vrE�a�ܮ�����  ��!���21��`( AAVM� �2�0 �@fd� TUP him� (J545� l)�`8 616� %�VCAM� ��CLIO] (�0:�5& � (F\ MSC ��Rt"PBsSTsYL�D!28 :2�\ NRE F2h S�CH6pDC�SU tpsh ORSR �r�D!04�SEI�OC& \fxh 542 LEX"� ESETn�8!H ���sh8 7H �OMASK�Ø"7>�.�OCO*`x�!0�3"6�!/400:66�$ G639.6[8LC�H!6OPLGR70=3
5MHCR��0�C� (! �06�A.�f8!54
��00D;SWb 588�180� �h!37 88 K(D�"02C24��N�27 q9�25���2-6�05��9�PRST bB/FRDMES�!zB��930 _ N�BA  6� HL�B 3 (~!SMވ@ Con� SPgVC �8!20z���TCP ara�m\TMIL� A��@PACET�PTX �@p T?ELN 96��2�9�%UECK��r� UFRM et��P!OR ORP I{PL%CSXC�0�j�1CVVF l� FQHTTP �stA")�I#� CG�HP8ZIGU�I�0�hPPGS oTool� H8�@�djZ��!@�h!6�3�%�@32Q\�31� B�h!96�%R6�51�Rs�!53 oTFAD�R41��8"1 ��oo�"9:��41775�"/@�P�VCTO�@�U�!�sh!80�%PRXyY�R�!770 �b~8 885 ol3P2� L� аdi� �`�ڳh LCP{Q� T'SS �b�26:���^�@CPE �HT@�VRC~�tQNLy ��@002 %�b	0dis� �`7� <��a\0�T�`1 ��`en�b4 6582�`)FU02Q0Π�o`p�Ptu�r4 d$r5N��RU0p@�nse�QJp1 A�PFI[ Jp3�g3}4�g40 al�xrE1t44w466� ts U0  7v��0O��r5�e�p7 �p "sw�a61d:��r4��r5 Qp!wGr`�$�p8R�"s�P`tQ�b�36w717�w8`�v83���r�8�&:��pOq8�8 _"rkey8�9F�v�a90�91 p�p#@��� �D095�g[97*pur�A1@ d���P|P�q1�0QplSq1p#4��]a!sM1@sl༂8��H��\1�d1�`��v��@{�14p�ae��5# h2��`�6ޣ��7�f1p@��d�YpCq(d�ـd�1�`uq���� Cu1< Oq� ��7&ReU1$ �u1�Pϱ�� ��@- WQ1�58 ase C渒9 B��60 �82ń�p���4 (Wai��`吢!���7E��8�EU1&P`ro9�<�1��<�2��<�	0��T��"l�5J�l��cC���9%�MCR��P��2�`�Q2@96I7�Q��8��9Z�A2TPB���P�2P7�U5@�o���
�58�`U���3 w����?A�E�1��c�qAw�l��A�1��512# f��1�u5Р��"�a5p$��56�+aĈ�Q5h��Ұ�1 �@��pp�b[�538 xaB��|p�4Ⱅ2�11/q5�p�4U=5�P16 (߲�P z��0��8�P��H���p�e5`�e5(�/�P`bbf>�X��$�Z�U�5d�\�� X�7 	  ~��8 k_kv���79 s�82 &�H5��E6���p�����h���ñ���3�J"�`��4 3Ȥ5�9ѧ6�0t���8Ⲗ6D0$�$�4 7���!���<�j67?0\tchk<�P`s��<�B<�90���7�<���<�\K�<�q �Ӻ�A�C<���q�<д��<�t��sg<�lIc���FA<�H���<���<Я���<�hk ��<Щ�B<е�o�<����<��K�<�dflar��<Ш��� ��@o�`���D�;�<�gEvam����B<гoќ���<а�KЀ�creexl����P�`��<���|���j6<�=s��prs.`��� \���<�7������fsgn��P�b�t�at��<�L��1|B !�svsch/ � �Servo S΋�ule>�SVS��44�1u�_<���� (����ched��,��~��A\�� �� B���B�qA�h���cj�� � 5�1<���Ә�p��css "ACS <�&(��6� ������c el���Q�����torchm�s�<�- T�Ma�`Ѵ���09 J5�;598 J681s�7� 8��b���<Чa����te,s�����/�E��� m��ARC..�� 1q�4�!=�,�C�tc�pA�@t����f� F����7#�2x�SE�r����UtmS�09610'���RC�������� p��96`G= '��"H5W�@���L���\f� � �PATb���`!a4U�#!Stmt��E ��� �pM�A�!p��z�2?�i�n_<�X��r�X e/cW����V����etdl�vߏ\oveto���܏���mmonitr`�\��|#�0st��?.6a��PP�����! Q�!y`�`asme �Arol�6c�43�0 �pl���01� 25��  �<� v	�v	�A>@�818\n; <�s�I�B�2�pMPT�P"��C�1mocol��,��CT�v�'!`� �A���8P53��y`Touchs�s0�`��<��J5��@�Ѩ`mP����n[P Q�a,�E�a��IPL&
�Pth�A<�KF#xR�m;�Qetth�THSR'�q-�Rt���o "PGIO��#!$s�ISwka�"cWK��!�MHqWH54��5w5n/"�Sm/��@ 7�*�da��8`!w/Ac��tsnf Tk�/�#@gb�a��u`��^m�`Au��Zӭ�ܱQp��@��#���Ka<��M��t5QtZ�a<��d�FS5GK����G�1o1r��dW��64��tP@x���P ����x,� �?$���P<�Z4e�7�g "SVGN�.ox�copy "CO;�Wj$�O�A�9� "FSG�ѧ�%�7��_��f� wQS�WF*!"(�sgat�uɀ���_
��tpN_TPDo��9�79�#dߎ?���h��GAT���!#��  �Гf�` �@�"/� �w�Z� �b?6 ?� ����� ���E �8��M� �chrT� �K6K� �sms� �o6��ѐ�gtdmen�?3 �?��� ���mkpdtd2 ���, ���pdQ�X� ������ ���mvbkup�. �[�C�С��mk3uno��prp���Gmkl �4��s ��niU��� �ldv9rw���glg�4��� ��棑��aut7�.pб�旐 �ַ������su3� ��@�� �Ƿ� ���\ �6�b2X� ��&�� �x����A4�  ���B   946�" ��fB� �t\p�aic\p4k947 ���F#���� ��ictas���pa`���cc:�<��8o�����gen�� �I ��F�lnp � �Ď��stf@��1��wbO�c��Ջ�`��߄�vri�ߢ�а�-T� ���p�flo�w� OPAc��ow���R50qtS �#T� (A��4�#�0��pѣV�cu3�Q0F� ��SI�ac�����46����s&��p�a��!!���� ���55�b �o)�p���0�|��
�afcal3�P� ��f��}���`�f��m	߳�p�d�m�/���a/��$C`ѷ��� �! trac�k\P� 0�ine/Rail Tr��]TJ�69W�T  (L��8(`љT.�`� %��D��P0� (��8�48��_ɛ�₇�4����� �3b�b3���alV@ �NTf���%��I�in]0m���aen������&?5�8c@Itst3@�� $����`�,R9�%����0氱%��po�peners-OW dDev��F�M�6W���|A�Pc"�l!esv� �,��R�V$�Q���U<�V$ �k)9j �6��# ��ȼ��%paop/!O�PNU�V ��2c#elL��8g_��8/�6��tscG��$Ѐ�V!�3� 5vrCop�ߡ�7`�n( `�V"2D�a V'O$�:S9��� Pump E��jQ�@�" ��!
��@бMSC#�@��)P���AC�`��� � �v���� \mh/plug�@g�"�7P��uK")㠱io�7�CJ0��E�LI�O q1g 7A93շ�5 q9 t����]4rb ST��R�ÞCPJ989�P�L�SE�' �e C3Q(P �/Ov���o�P� ? I1�R����55��f�I1`�tcwmio��MIO������Utco1"CL�01V �cBK`iEo��uM?���Sl� I0�ߢ�Eg �o���fb �tI4\onfdtI����e%�p27�Inste�TB CoMIoo1E�R�(do554 (;r>Ex�,��nR##ipc��/>��qp5���
@oQé�1�p����7/o����ra�pd�CD V_��rP�֮��qp2Gcnd��s �p��a�o�r`҄�S��"�bc�a�c���2kI�<�?A�pcrt���or0�qd#��"���3p�+���D��Џ��vr2k�0���AG�.�+��cho�;�u�C��(� �uV630 �fwe P�mී�@�X��`��TX�� ��>d�chp "_��(	�3�����8����\p3�v�������9�3�1 ������low�[ͧ���c!hk���㳦s��s?Ө0�i�1h���2�� i�w����s?1*�`-	�:�O��vr�������0�'���PFR�APWat?1rn�eE�P�sp�& ac5�� _A�rbo#�, �a��g�������z�Qs<�ICSP+� 9_����� ��F�A9PH51�IQ93 7��HX6�hQ]PVR`S5��fPR�6 iQWPR� (�P!am S�u�"�A�I0�tppr�g�0���`h�@2atk932�!��E��^��asc "8�C8��S>i�atp�"��d�@1I�
g�ds�blfltJA�Qs�able Fau�P{C!��EV0ex~/!DSB (DC��t�$�p��X 7�@� �� 5��Q�t3*��~���td9� "`!%�(5��sb9������\	�6#���@�5�p$D@550-A�djust Po'intO"tVJ�Rs�z�䐄��!�X_�Yj���0\sg��4x��}7y�\ada�O"ADJ���j�Q�etsha<�SH�AP�sŭ'jpo �r4�t�!��$ �(�C|�	Tk!bRP�KAR/Qiagn/ostì!O!vV66 J`ew0��(�L���/�&krlde� ��PP�� �hU b���r3�Pyp?q��DBG2C��� �X�o�1U��� ��WT`�@i�pJCM�aipper Opv`1Se}�78 (MH G F� ;":�&##�� a��x�֕$��388�C�����#��9.�9�C��g##PPk�Q��8 �!�_"$�"��=0%�P� �A $��_�#%0AQ�C�~2 Mat.HandlE��!= &�pq MPLGET�0�1(�3�Tt&P�Sٰ' �B�1��B0����&p� �H��PP �'p��@�C 7PP	�TG�tD5�}�m�q�Afhnd �"F_R  ������PP	   pxT?Q���P(Pa���To�����?�p�mpaO��JP ak925��2`@O�JR	psQ`B2�unLHP�T7gse�GSo1�O�W�QT��v !�R��Ptp~���JRdm�on.�@��V�!ns�hYvr�QJ�g�Q`�o�jY�HS~7sl�f] ��pen�PDnRp(R&���ɐ823'� �ٔq���g� ����� 1�� S�� ? �c\sltQ�!|QE�P��a �rtPg��P�� �v��"SEDG8�s0.�qtdgY T�� ��vP`ho�s`<` ����qc�`g
�e`� o�w�a@o"�ile6�H�e�ȅnR��� �e! j517�>Ճ��J%��e�`��Q4��Q&�!L�!F�J�=�o�5�z/l17���_�œ���`C0C�  ���LA/NG j��A��p������gad����#�jp�.`��4�Ē�ib�0��s�Ƒpa����&���j539.�f�,Ru� Env
�����2�3H�z�J9������h�Ф
Ҕ���2��2���� (K>L�n-TimФ������p�3�TS�����\kl�UTIL�"o���x�r "QMGl��!������1 "��S�T3�\kcmno��SФ�T2���ut�.�l�readc�}�exPY�ܤ�r��\��l�҄Фw�3��2C�*� -�C�D�E!Ĥ� .�4�C� R CV̴�҆��\p�Р���p�tbox��.�@��cycsL�:�RB�TE�veriOPTNE���;ӕӂk�e�ߦ�a�ߦ�h�g�ߥ�DPN��g�p.v��r�ptlit��0�4��te\cy���>�tmnu3`�r�����5UPDT�������駣���ite �� sw�to�,���oolB�F"�Y���Q��(q��gr3��䪒���"�䴁w������߳��s��������������lS���bx A"O�� ����l��`��P���A�l\t��� ��������	�Co�l�e!��R C ��r��&r �m;`��Chang�Lq�T1 �rcm3�"��
� 6���"����sPa7���"��22B2��2D4�57�� CC�FM�H��accda��Q�c' ��KÕ0���K!����m o!���,$Á��! "
����/�/����	�Y�,$��)�,$sk(����m rC%tS1,$�+��k1�%unc.�,$oñ�1��sub������1��cce �5/!&��-/?-W/i&vs�}/�%#�#�/��.C��/� C%
�@?  U �&+��F:qt�
pD�Ѓ D	 � U�:7�Dxmov.�P��DPvc\5Q�tfr@PeC_~UYgeobdtg_y[tu���P���PTUIt�P�Sx�_�^z�_��\var�_�\xy\�_�[pcl`c�P脆�P�Ue�Pgri�psuaoskuti����ovfinfpo}��o�j�b�P���Qud\�aX��Pc�\Rrp�Qnƅ�P�v�P)t�m#qƆ�P�v�a+ro�g�a��\Q�?a+rp#al?a{�{spa��@�P�u�Q�t�_TZp�0<�osipkag3r�o>vlclay(�:�t�pT�d�pu?a�c�A������KtKa�P䒏��qTf|rdm��{rin#r���As� �2���|s�PLd�v�tv��v�h�0��ystn* џ�y%t'�1�p��D�p�uϑ#�ul�@o�W6�92�siupdl�]�Fo�vr�on��`1L��z�`\�r���il3�$|l4��ǉ#q5 4FyB�Տg{�`���{�wcmס���wxf�er�UYtlk2�pp߿UYconv��sicnv�Qʯx�ag��H�Z�lct�`ao�=�p��׭nit0믁�3�������  �� ?v	�v	$��alϑpm�r&�B�eWa���f�%�� ����I��߬�u�ͬ�KamT�f���c��w��roǁ#�5�����?� sm��y�a��y� ��������`����͐ϑ��p��m�Wa� 1���A�6�S�e�X� �ψ�\Q}��������� ��ĥw߉�西߭�� �߮�#q0��rs�ew����1�a��z긱n�@�.�۲;�d�������  � �Ad	T$�1 �p! P��e �Ne 	lf@C��@�s/�  ?�����8�� �������r�eg.�C=��o�99 ~@�����$FEAT_�INDEX  �z ���e� ILECO�MP :��=�1!!z�$#SETUP2 �;1%;"��  N f!$#_A�P2BCK 1<~1)  �)��/�/  %�/�/e4 �/�/>%�/$?�/ H?�/U?~??�?1?�? �?g?�?�? O2O�?VO �?zO�OO�O?O�OcO �O
_�O._�OR_d_�O �__�_�_M_�_q_o o�_<o�_`o�_mo�o %o�oIo�o�oo�o 8J�on�o��3 �W�{�"��F� �j�|����/�ď֏ e������0���T�� x������=�ҟa��� ���,���P�b�񟆯 �����K��o���� �:�ɯ^�����#� ��G�ܿ�}�ϡ�6� H�׿l�����ϝ���t@)t Px/ 2� *.VR��߅�*�@߂�F�j�T���PCrߛ߅�F'R6:����V���z�T �!���K�� ��q�S�*.F�ߢ��	�Ӑ���x^����STM ��'���S����iPendant? PanelS���HI���9���U�������GIF0;�p�������JPG���;��]oR�
�ARGNAME.SDTy�>�\"����Rc	P�ANEL1Y�%�>��e�w��2 �A/�//���/�3_/�/��/p/�/?�4�/I?�7?�/?��?TPEINS�.XML�?>:\��?t?�1Custo�m Toolba�r�?Q�PASS�WORDg?w�F�RS:\:O�? %�Passwor�d Config {OR��OSO�O�O��_ �OB_T_�Ox__�_�_ =_�_a_�_�_�_,o�_ Po�_Io�oo�o9o�o �ooo�o(:�o^ �o�#�G�k ���6��Z�l�� �����ƏU��y�� ����D�ӏh���a��� -�Q��������� @�R��v����)�;� Я_������*���N� ݯr������7�̿޿ m�ϑ�&ϵ�ǿ\�� ���y϶�E���i��� ߟ�4���X�j��ώ� ߲�A�S���w��� �B���f��ߊ��+� ��O���������>� ����t����'����� ]�����(��L�� p��5�Yk  �$�Z�~ ��C�g�/ �2/�V/���// �/?/�/�/u/
?�/.? @?�/d?�/�?�?)?�? M?�?q?�?O�?<O�? 5OrOO�O%O�O�O[O �OO_&_�OJ_�On_ �O_�_3_�_W_�_�_ �_"o�_FoXo�_|oo��o�o�`�$FIL�E_DGBCK �1<���`��� ( ��)
SUMMA�RY.DG�obl�MD:�o*n`�Diag Sum�mary+8j
C?ONSLOG �qn�=qCon�sole log��7kpMEMCHECK��2���qMemory� Data3�;g�� {)�HAD�OW(�����C��Shadow C?hanges���c�-��)	FTAP�����=��q�mment TB�D;�;g0<�)�ETHERNET�0�`n�q~���=qE�thernet ��pfigurat�ion��B`%�DCSVRF/��'�@��C�%� ve�rify all�C��c1p� �DIFF8��0�ůD��%Z�diffǯ{��q�1�������J� X�q�|�=	�CHGD�&�8�ͿD�ܯ������2Ŀ����R� `�yτ�GD�.�@����D�����FY�3�ϳ���Z� hρߌ�GD$�6�H����D�����UPDATES.$��
�ckFRS:\�"�c�>qUpda�tes List�c�`{PSRBWLOD.CM��blN����e��pPS_ROBOWEL\�6o+� =�loa��o����&��� J���n�����9�� Jo���"��X �|#�G�k �d�0�T�� �/�C/U/�y// �/�/>/�/b/�/�/�/ -?�/Q?�/b?�??�? :?�?�?p?O�?)O;O �?_O�?�OO|O�OHO �OlO�O_�O7_�O[_ m_�O�_ _�_�_V_�_ z_o�_oEo�_io�_ zo�o.o�oRo�o�o�o �oAS�ow� *��`���+� �O��s������8� ͏ߏn����'��� � ]�쏁������F�۟ j������5�ğY�k� �������B����x������C�үg�v���$FILE_N�P�R]���Y�������M�DONLY 1<���U� 
 � �ۿ(���L��5��� Y��}Ϗ�ϳ�B��� ��x�ߜ�1�C���g� �ϋ�ߘ���P���t� 	���?���c�u�� ��(����^����� ��$�M���q� ����� 6���Z�����%�� I[���2�����VISBCK�����ų*.VD��*� FR:\�V� Vis�ion VD fileVd��� ����	/./�R/ �v/�//�/;/�/_/ q/?�/*?<?�/`?�/ �??�?�?I?�?m?O O�?8O�?\O�?�?�O !O�O�O�O�O{O_�O !_F_�Oj_�O�_�_/_��_S_�_w_�_o~�M�R_GRP 1=LeC4 w B�`	 ���lo~li`۬B���D��f�nӺMT� ��� ����e `i`a�o�khb�h�o�d�cic.N��BL&�2L��N��dH��E��|��i`?5�
A�O�@
\=>�aA�88���l}A�A�ڛA�}�s����p�l}F@ ��qhq�y�~g�fF�6�D�MqD��� BT��@���Ô~pD��6����l���5��5��|���~�?B�C��Bpm.Bx��A�akBWqr��~T8�B)+�B4�A���aB#�`l叐�A�����A�܏�e�P���t�����@�bo=���@�	Ƙ����Ο ��+��O�:�_���`p�����eBH`� �����a?�ŉ��'�d
���Z��WZ��a�/�FX
�A@�~��@�33@���'�\��[���ѿ��@��񿋯�*���N�9�r�]ϖρ�<��G�=�<��m]<�+=~��m<c^��8�eN7��7�ѷ7�x7;��51���	ߤϨ�?߾d2^`Yb`�*b`�����F�`�U�b` b`�0�����C�^o�߂o�o �߸o��o�� ]�(� ��l���������� ��#��G�2�k�V�{� �������������� 1 ��-�) �������0 T?xc��� ����/')�'/ M/_/q/8��/�//�/ �/�/�/?#?
?G?2? k?V?�?z?�?�?�?�? �?O�?1OOUO@ORO �OvO�O�O�O�O��_ ��J����`_*�_N� �_�O�_�_�_�_oo 'oMo8oqo\o�o�o�o �o�o�o�o�o7" [Fjh�x� t��!��E�0�B� {�f�����Ï���ҏ ����A�,�e�,/�� �������/�J��� �=�$�a�H�Z����� ����߯ʯ���9� $�]�H���l�����ɿ ��ƿ���#��O�OV�  _z�D_V_��z_�Ϟ_ ���
�C�.�g�R� ��vߛ��߬�����	� ��-��Q�<�N��r� ���������)� �M�8�q�\������� ����������7" [Fk�|�|�� ��֟3�WB g�t����� /�///S/>/w/b/ �/�/�/�/�/�/�/? ?=?(?:?s?:�LϦ? p��?�Ϧ� O��$O�� T?]OHOZO�O~O�O�O �O�O�O�O_5_ _Y_ D_}_h_�_�_�_�_�_ �_�_o��@o
�go*o wo�o�o�o�o�o�o	 �o-*cN�r �������)� ;�M��������� ˏݏď��%��I� 4�F��j�����ǟ�� �֟��!��E�0�i� T���x���ï�?�?�� O��?OO�t�>O ������ѿ��ο�� +��O�:�s�^σϩ� ���ϸ������ �9� $�6�o�6o��Zo��R� ���������5� �Y� D�}�h�������� �����
�C�U��y� ����d�����:����� +Q8u`� ������ ;&_Jo��� ���//گ4/�� x�j/4��/X�n/|��/ ��/�/!??E?0?B? {?f?�?�?�?�?�?�? �?OOAO,OeOPO�O tO�O�O���O�O_�O +__O_:___�_p_�_ �_�_�_�_�_o oo Ko6oooZo�oZ��o�o �o�o��xo
G2 kR������ ���1��.�g�R� ��v�����ӏ���	� �-��Q�/*/��N/ ��r/�/ޟ�/��/)� D�M�8�q�\������� �����گ���7�"� [�F�k���|�����ٿ Ŀ���O�O�O��W�B� {�fϟϊ��Ϯ����� ����A�,�e�P߉� t߆߿ߪ��ߪo�� +�=�a��߅�p�� ���������� �9� $�]�H���l������� ��������#G2�W}h�p��$F�NO ������W
F0� �  #��1 D|�� R�M_CHKTYP�  � �q�� k�� ��OM� �_MIN� m���}�  X� �SSB_CFG �>� ~�Jl�Aj|��TP_DEF__OW  m��>�IRCOM� ���$GENOVRoD_DO���n�THR d��d�_ENB� ��RAVC_G�RP 1?3� X�e/��/�/�/ �/�/�/�/�/? ?=? $?6?s?Z?�?~?�?�? �?�?�?O'OOKO2O oO�OhO�O�O�O�O�O\�O�ROU? E�. q����>��8�?#�O_�_K_m_o_ꐖ  D3���_E�_q�@A��\Bȡ��R���>Y_6 SMT<#F�C-�Ufoxo�o�HoOSTC,1GYn?��_ 	�hM�k�o�f�oyeCUgy �z1�������p	anonymous�5�G�Y�k� w��o�o�o���� ��*�<��`�r��� ����ˏ	����� &�8������������� �ȯگ���M��4� F�X�j�����ݟ��Ŀ ֿ���I�[�m�ρ� fϵ��ϜϮ�����}� ����,�O�Pߟ�t� �ߘߪ߼���/�A� C�(�w�L�^�p��� �ϸ����������a� 6�H�Z�l�~������� ����9� 2D V��z������ #��
.@���� ����������� //g</N/`/r/�/ ����/�/�/?Q cu��/[?��?�? �?�?�?)/�?O"O4O FOi?�/�/�O�O�O�O�9m�aENT 1H�[ P!^O_  `_?_._c_ &_�_J_�_n_�_�_�_ o�_)o�_Mooqo4o �oXojo�o�o�o�o �o7�om0�T �x�����3� �W��{�>���b��� Տ���������A�� e�(�:���^���������QUICC0 �̟ޟ?��1@��.����2��l�~�߯�!ROUTER�௼�ί/�!PC�JOG0��!�192.168.�0.10	��GNA�ME !�J!�ROBOT���NS_CFG 1G�I� �A�uto-star�ted/4FTP:?�Q?SOBχ?f� xϊϜϮ��?������ �+�߿�P�b�t߆� ��6�����(�J�  �1�C�U�g�6ߋ�� ��������x�	��-� ?�Q�c� ?2?D?���� �����)��M _q����:�� �%t�����m ��������� �!/3/E/W/z{// �/�/�/�/�/6HZ  ?n/S?�w?�?�?�? �?�/�?�?OO<?=O �?aOsO�O�O�O�/
? ?.?0O_d?9_K_]_ o_�_PO�_�_�_�_�O �_�_#o5oGoYoko�O �O�O�O�_�o&_�o 1Cogy�� ��oT��	��-� |o�o�o�o����o�� Ϗ����)�;�M� _�q��������˟ݟ��ÿT_ERR �I�����PDU�SIZ  �^ڴ��$�>=�WR�D ?޵w�� � guest+�}�������ů�ׯ��SCD_GR�OUP 2J�� �`�1��!怒L_���  ���!�	 i-	��E���Q�E� EATSWIL�IBk�+��ST 4�@���1��L�FRS:�аTTP_AUT�H 1K�<!iPendan�������!K?AREL:*���	�KC�.�@���VISION �SET���u���! �ϣ��������	�߀P�'�9߆�]�o޽�C�TRL L���؃�
��F�FF9E3��u����DEFAULT���FANUC� Web Server��
��e�w� ��j�|��������WR_CONFI�G MY��X����IDL_�CPU_PC�惑B�x�6��BH��MIN'��;�GNR_IO�K����"��NPT_SI�M_DOl�v�T�PMODNTOL�l� ��_PRTY���6��OLNK 1N�ذ�� �2DVh��MASKTEk�s�w�Oñ�O_CFG��	U�O����CYCL�E���_ASG� 1O��ձ
  j+=Oas�� �����//r.�NUMJ� �J�� IPCH�x��RTRY_CN��n� ��SCRN_�UPDJ����$� �� �P�A��/����$J23_�DSP_EN~���p�� OBPROqC�#���	JOG��1Q� @��d?8�?� +S?� /?)3POSRE�?y�KANJI_B� Kl��3��#R������5�?�5CL_�LF�;"^/�0EYL_OGGIN� q���K1$��$LA�NGUAGE ,X�6�� vA��LG�"S�߀���J��x��i��@<𭬄�'0u8������MC:\RS?CH\00\��S@�N_DISP �T�t�w�K�I��L�OC��-�DzU�A�zCOGBOOK U	L0��d���d�d��PXY�_�_�_�_�_ nmh%i��	kU�Yr�Uhozo�hS_BUFF 1-V��|o2s��o �R���oq��o�o# ,YPb���� ������(�U���D/0DCS X>u] =���"lao�����ˏݏ�3n�I�O 1Y	 �/,����,�<�N�`� t���������̟ޟ� ��&�8�L�\�n���@������ȯܯ�Ee�_TM  [d� (�:�L�^�p������� ��ʿܿ� ��$�6� H�Z�l�~ϐϢύd��SEV� ]�TYP�$���)��m�1RSK�!O�c�"�FL 1Z�� ����߯���������L	�:�TP5@���}A]NGNAM�$��E��k�UPS PG�I|%�1�%x�_L�OAD0G %Z%TEQѼ���MAXUALRM ;'�I(��~���#� QV�#a��CQ[x�@8��n��"�1060\	 �F�	�Ϣ��� ���������� D '9ze���� ����R= va������ ��*//N/9/r/�/ g/�/�/�/�/�/?�/ &??J?\???�?k?�? �?�?�?�?�?�?"O4O OXOCO|O_OqO�O�O �O�O�O_�O0__T_ 7_I_�_u_�_�_�_�_��_o�_,o��D_L?DXDISAc����MEMO_AP�]�E ?��
 �5i�o�o�o�o��o�o�o��ISCw 1]�� �o Td��\no�� �������I� 4�m��f���$����� ����!��E�ƏT� f�:�����ß����� z��ܟA�,�e�w�^� �����~������  �=���L�^�2����� ����߿�r� �Կ9��$�]�o�(t_MST�R ^�͂�SC/D 1_xm�W��� S�������=�(�:� s�^ߗ߂߻ߦ����� ��� �9�$�]�H�� l������������ #��G�2�W�}�h��� ������������
 C.gR�v�� ���	�-Q <u`r���� ��//'/M/8/q/�\/�/�/�/�/�/s�MKCFG `����/��LTARMu_2a��2� �#\`Y>G`M�ETPUT`�"�����NDSP_CMNTs506�5��' b���>�"1��?�4�5POSCFz�7�>PRPM�?��8PSTOL 1�c2}4@p<#�
aA�!aEqOG]OO �O�O�O�O�O_�O�O A_#_5_w_Y_k_�_�_�_�_�Q�1SING_CHK  +O�$MODAQ73d�
?�7:eDEV �	��	MC:>MlHSIZEs0����eTASK �%��%$1234?56789 �o�e�gTRIG 1en�� l��%��?   A$�Üf�YP�a,u��cE�M_INF 1f�>7 `�)AT&FV0�E0N�})�qE�0V1&A3&B�1&D2&S0&�C1S0=�})GATZ�� �H� E��q9m��xAu��� X�������� �� ����v�)���я ��П�������*�� N�����7�I�[�̯ ן���9�&���\� ���g�����i�ڿ�� ����ï4��XϏ�i� ��A���m�������� ��ѿB����ϊߜ� O������ߟߩ���� >�%�b�t�'ߘ�K�]� o߁�����(�_�L� ��p�+����������.�ONITOR�0G� ?ak   	?EXEC1�#U2345T�`789�#��xxx *x6xBxNx@Zxfxrx2U2�2�2�2�U2�2�2�2�U2�33�3�aR_GRP_SOV 1g�y�a(�Q�>`^�?������žee@?�<I�����Ƥa_Di�n�!PL�_NAME !��5
 �!De�fault Pe�rsonalit�y (from �FD) �$RR2�� 1h)deX�)dh�
!�1X d�/d/v/�/�/�/�/ �/�/�/??*?<?N? `?r?�?�?�?�?�?�82S/�?O O2ODOVO hOzO�O�Ob<�?�O �O�O�O_"_4_F_X_�j_|_�_LhR� 1�m)9`\b0 Ә_pb�Q @oD�  �Q?��S��Q?`�QaAI�Ez  a@og�;�	l�R	 '0`4b@4c.a��P�Jd�Jd�K�i�K�J����J��J�?4�J~��jEa�o-a�@��o�l[`�@�z�b�f�@�S��a�Q�o�c��=�N��
������T;f���`��l[`�*�  �p  ��$p> p�$p��o?�p?����������o�B ntr�Q�skse�}�l��p�  |�pu`j  #p���vks�� 	'� � ��I� �  ����}:�È~6�È=���N��b@^�d��n�Q����{�R�x���nN<. ��  '���a��`@a�@�t��@p@p@-CpC0�f0�+p�B/pC3}�P��@%�Eab��oo$|m�/���gA%���. ���z�`�P���QDe���˟��(���m�� �t� O� ru� �4 �xR�c��s� :	e�a�P�` �?��ffb�!�����7� ��گ쬛af���>搠���iP��P;�e�S�Ea4f�u��>LX��s�b<	��I<g�<#��
<2��<D?��<��
vo���¯�S��S.���?offf?u�?&�ޗd@T���?��`?Uȩ?X����Z���T:z �TB��Wa�з*dů�� �Ϻϥ��������&�`8�#�\�h�+�F.  Kߘ�G߼�3���Wɯ����G�@ G����X�C�|�g�y� ���������jZ�� �ￏQ����ߙ��� ��3�������/ A��t_�����������b�� �@+Fp�IP(�t��%���[`B�0����<ze�cb!@I��
�M`B@���@`�9@y���?�h� ��@�3�[N���N�N�E��<��/:/L �>���ڟ�A�p��C�F@�S��b/DpX������@�t��%��h��`/qG���GknF&��FצpE,8�{�/ F�Z�G���F�n�E�DE,ڏ��/� ���G���F7��F��ED��.��C?.? g?R?d?�?�?�?�?�? �?	O�?O?O*OcONO �OrO�O�O�O�O�O_ �O)__M_8_q_\_�_ �_�_�_�_�_�_o�_ 7o"o4omoXo�o|o�o �o�o�o�o�o3 WB{f���� �����A�,�Q� w�b����������Ώ ���=�(�a�L����p�����(r!3�j�i��r���ꕢ�3�Ա�ڟ�u�4 ����u�Pq�2�D�&�jb^��p�1w���������ʯ���ܯ�� �s�P^�PD�c� `�m���y�\������Ӱ�¿Կ����� .�G����}ϳϡ� ��홍�U�_�J���$�y.�@�v�d�z߈� ��x�4�������� �h�D�.�2� �$[�'G�[�^�B���B��CH� ^�� ��u�����������p�h�M�_�q�����T�����^�^��Y�m�2��
  ����#5GYk }������h*��� ��>�x}���$MSKCF�MAP  ��?� �����m�N"ONREL7  6�9_��"EXCFENB�k
7]�FNC��}JOGOVLKIMkduyd"WKEYk�"WRUN��"SFSPDTYU�x�v_SIGNk>}T1MOT�z�"_CE_GRoP 1n��9\���/���/�/4��/ ?�/2?�/'?h??�? C?�?�?y?�?�?�?O �?@ORO	OvO-OoO�O cO�O�O�O_�O*_<_�#_`_-�"TCOM_CFG 1o/����_�_�_
|Q_/ARC_�6��UAP_CPL�_��NOCHECK� ?/  5�;h9oKo]ooo�o�o �o�o�o�o�o�o#�5GTNO_WA�IT_LF'5y"NMT�Qp/���qo_ERR�!2q/_�� R_����"�:�L�dT_�MO�sr�}, ��jP_��_�PAR�AM�rs/�������MW��� =�e�345678901.�@�R�)�q��� _�����˟����ݛLW�3�E�؏i�c�UM_RSPAC�E,�������$ODRDSP�SI&��OFFSET_C�ARToݨDIS��ݢPEN_FI�LE�I!�Q�v�PO�PTION_IO����PWORK kt�'� T�|�
�@^�F�U��Z���	 �m���C��
���RG_DS�BL  ��v����ޡRIENTkTOj�C����8�ῠUT_SIM_DJ�6	���VàLCT u��}\��Q��W�_P�EXE���RAT����� ���UP� ve������`�����*�8��$���2�#h)deX)�dh�O�X dY�ߑߣߵ����� �����!�3�E�W�i� {������������2n��)�;�M�_�q� ��������<��� ��+=Oas@���X��� O���1m(���(��.�g��"0 �дu�  @D7�  �?���?рH�D4  �EzZ3;�	�l	 0DӀS@SM� �i��i �H)!H�,�H8�H�m�G�	{Gǎ8��6�MV���� �C�)����)����Ճ�*�  �p  �
 > � ,�//�)/ B,�Btr߰«�H�¼�/���/�"`�# �,0 �� _�  � ߽poj  B ��&�X�?MU	'� �� 12I� ��  ���-=����U?g;/�@}?�0~.ѱ�?;Ѳ����H[N5��? � 'M�D�> C)�f)�J BN +��=x%O7O�R�@D1~�oo$�����JWA�D0�J5�4�:  �1�E&?�O�O#_�_G_2]�� ��t O� �ru �4 ���R�Uɳ� :��%S�р� �?�ff��@[�_�_BV_{�o~��18р�"o0j>�P�Q6YP�рZo�WrAdS�%��>Lw0�#�<	��I<g�<#��
<2��<D��<�ל���_��j�ѳMb�@?offf?�0?&p�:T@T�q?��`?Uȩ?X�-q�iyBq5Y a��gI�_� �����!��E� W�B�{���d�����Տ�LnpΏ/�ʈG�@ G��U�ȏy� d�������ӟ����� ��yB=� ��?p�� �/򏸯�߯R��� '�9��oN�`�����~�P����ۿƿ�B�� �D�e�ֿ;�ҿ_�J�?��h�oϨϓ�J���D4��b!�_@ ���� ߧ��Ŀ�����%�@I�)�M`�B@��@`��9@y��?��h	� �@�3��[N��N�N��E��<�/�Y�kЖ>��ڟ��A�p�C��F@�S���pX������@��t��%�h���߉!G��G�knF&�F׿�pE,8{�� �F�ZG����F�nE��DE,ڏ������G��F7���F��ED��Mf��b�M��q�� ����������(�� 8�^�I���m������� ��������$H3 lW�{���� ��2VAS �w������ /.//R/=/v/a/�/ �/�/�/�/�/�/?? <?'?`?K?p?�?�?�? �?�?�?O�?&OO#O \OGO�OkO�O�O�O�N=(]�3�ji�O�a���	U�E3Ա�x�O_<q4 ��%_<7_<q�P�Q_c_�ERjb}_�_1w?������]�Y��_�_o�_1ol��P�bPcn~���o�O@�o{_�o�oY�`��o �o,/;M#�f 0o�����Y�e@t�~�i#�1�C�yM� _�����������{bS� Ԏ��	�?�-�c�Mj�2���$�VG�Dz}�B����B��CH�}�9�֟��� ��0�B���wl�@~�������Ư�T�E��\��qQ��U
 ί�0�B� T�f�x���������ҿ����χ��� ���]{x}��$P�ARAM_MEN�U ?Յ��  �DEFPULSE��	WAITT�MOUTl�RC�V� SHE�LL_WRK.$�CUR_STYLvj���OPT��N��PTB����C��R_DECSNw� Te'�!�3�E�n�i�{� �߶߱������������F�A�USE_P�ROG %P�%�B��V�CCR���UeXÚ�_HOST7 !P�!����Tt`����������4���_TIME��� �T�  A�GDEBUG��P�V��GINP_FLM3SK]���TR����WPGA�� |�[����CH����TYPEM�Y�A�;�Q zu������ 
)RM_q �������/ */%/7/I/r/m//�/��/�/�/�/?��WO�RD ?	��	�RS��CPNeS�E��>2JO��ξBTE���TR?ACECTL�PՅ�Z� {`�/ a`{`�>�q6DT QxՅ��0�0D��Sc7{a�0����2���?�?�2��4D�2#A�O.O@ORFcA�bBU`D	`D
`D`DU`D`D`D`DU`D`D`DObOtO�F A�5P�2 Q0TOBPRPBP�BP0T�BP�BP�BP�A,_>Z�_=_ O_a_s^$_�_�_
b�� "o4d�_�_�_�O�O_P_a�1	ad�TUVd^dfdnb�Wr�k}�o�o��j;qwc�TvT ~T5OcM_q�� ���v,>�
�t �@�R�d�v������� ���6,�>�P�b�t� ��������Ο���u �9�*�<�N�`�r��� ������̯ޯ��� &�8�J�\�n������� ��ȿڿ����"�4� F�X�j�|ώϠϲ��� ��������0�B�T� f�xߊߜ߮������� ����,�>�P�b�t� ������������ �(�:�L�^�p����� ���������� $ 6�Fl~��� ���� 2D Vhz����� ��
//./@/R/d/ v/�/�/�/�/�/�/�/ ??*?<?N?`?r?�? �?�?�?�?�?�?OO &O8OJO\OnO�O�O�O �O�O�O�O�O_"_4_ F_X_j_|_�_�_�_�_ �_�_�_oo0oBoTo foxoN�o�o�o�o�o �o,>Pbt �������� �(�:�L�^�p����� ����ʏ܏� ��$� 6�H�Z�l�~������� Ɵ؟���� �2�D� V�h�z�������¯ԯ ���
��.�@�R�d� v���������п��� ��*�<�N�`�rτ��ϨϺ����$PG�TRACELEN�  ��  �_�������_UP y������������_CFG �z����� ���<���N�V�h�r�$�D�EFSPD {�/��������I�N'�TRL |�/���8Pի�PE�_CONFI+�}>���<�]x�LID(�~/���GRP 1���������@��
=�[���A�?C�C
�XC)��B��r������dL�z�������� 	 xr�Nߣ�  ´�����B������������A���> �6>7�D_�������� ='�=)���������	B -��Q�M����  Dz����
 ��&L7p[ ������/��6/!/Z/��
V�7.10beta�1<�� B=}q�"`ff@��"�>����!=�{�͏!A>ff�!�@�ff�"�\)��"D��?�  b�!@�!� �!Ap�#W��h/??*?<?K;#�w����O/�? K/�?�?�?�?O�?O >O)ObOMO�OqO�O�O �O�O�O_�O(__L_ 7_p_[_m_�_�_�_� �_ o�_$oo!oZoEo ~oio�o�o�o�o�o�o��o DQy{/�#F@ {yw}�y{� �y�-������/� Z?l?~?w���t����� я���������O� :�s�^���������ߟ �ܟ� �9�$�]�H� ��l�~����_ۯ�� ���5� �2�k�V��� z�����׿¿����� 1�\n�j�|϶� ������	�4�F�X� j�c�χߙ߄߽ߨ� �������)��&�_� J��n�������� ���%��I�4�m�X� ����ί���������� !E0B{f� �����H� Zό�Vh�ϴϊ� ���� �2�D�V�O/ �s/^/�/�/�/�/�/ �/�/? ?9?$?6?o? Z?�?~?�?�?�?�?�? O�?5O OYODO}O�O ���O�OtO�O�O_�O 1__U_@_R_�_v_�_ �_�_�_�_"4Fx Bo|����o��o �o//0/B/;�__ J�n����� ��%��I�4�F�� j�����Ǐ���֏� !��E�0�i��O^��� N�ß՟������� A�,�e�P�b������� ���o o2oTo.�ho zo�o�����o��Ϳ�o 
گ'�֯K�6�o� Zϓ�~Ϸ��ϴ����� ���5� �Y�D�Vߏ� z߳ߞ���������� 1��Uy��:�� ��������	���-�� Q�<�u�`�r������� ����T�f�x� n��������� ���7"[F j������� !//E/0/i/T/f/�/ �/�/�/�/�/?�//? A?l�e?w?&?�?�?�? �?�?�?�?OO=O(O aOLO�OpO�O�O���� *�O_@RdZ_l_���$PLID_�KNOW_M  ���|�A�TSV ����P� [?�_�_o�O&oo#o�\o�B��SM_GROP 1��Z� dI`��oo$�Cf�d����D��TPbj�oLk�f �o"~�U�o>n 2T�~���� �7�4���p�D��� R���ʏ���������� 6�
�T��*������Q+MR�c��mT�EGQK? GR��(�#� ��[��/�A�S����� �������$����W� �+�=�O��������� ��� ���S�Ͻ�{ST�a1 1�������P0� @����E�ϲ����� ����M�0�B�T�f� �ߊߜ����������ߠ7��,�m��2������A�<��z�3 �������4���������5)�;�M�_����6x���������7 ����������8(�:L��MAD  ����� ��PARNUM  ��qKo���SCH�
 �
��S+UPD��xaq{>��_CMP_�`� �<Pz '�U�ER�_CHK���0�Z���RS���_��Q_MO� �%_���_RES_G
����� ��v/{/ �/�/�/�/�/�/�/*? ?N?A?r?e?w?J'��W,g/�?L%��?�? �?N#(��?OON#w� 4OSOXON#��sO�O�O N# �O�O�ON#d �Ox__N"V 1��U�ua�@cX��Pp��P$@cW،P���P@@cV��P��"THR_INR����pbA%d�VMA�SS�_ Z�WMN��_�SMON_QU?EUE ��e���`Ȩ`�N�U��N�V�2`END84a6/NiEXE]oNe�WBE\`>o/cOP�TIO;g?+2`PR�OGRAM %�j%1`O_�0bT�ASK_I��nO?CFG �o��9pDATAɓ�.B{@ev2w�� ����z��+�=� O��s���������nz�INFOɓ��}� !dr��!�3�E�W�i� {�������ß՟��� ��/�A�S�e�w�҇ބ��| �98q�?DIT �Bׯ>j~WERFL~hwS�~�RGADJ ��ƪA�  ,�?�E�8��Q�IORI�TY�W���MPGDSP�a�j�U�W�vT�OG��_T�G���Rj��TOE��P1�ƫ (!AF�PE5 ���?!tcp��%͟!ud�?�!�icm<�Q_��X�Y_<q�Ƭ�Oq)� *������Op���������� ��<�#�5�r�Yߖ�}߀���߳������&�*��PORT�a��OpA%�_CARTREP~`Ʈ���SKSTA�X!*S�SAV`�ƪ	�2500H809�u�T毙䕣�ƫ
�����`X#�$��6�m�URGEU`Bl��A)WFP�DO�V��2�W�q�?Q�W�RUP_DELA�Y �Ưe�R_'HOT�hwR%z�����R_NORMA�L�n��6SEM�I:y�QSKkIP���X%�x 	������ ��X%-;%[ mE����� ��!//E/W/i/// y/�/�/�/�/�/�/? �/?A?S?e?+?�?w? �?�?�?�?�?O�?+O�=OOO1U�$RBT�IF��NaRCVT�M�����m@DC�R����AA�.�B�{A��).?� �@���)�������c/ž�=B����[�_� <	�I<�g�<#�
<�2��<D��<��
+__{_�_)` ���_�_�_�_�_ oo $o6oHoZolo~oi_�o �o�o�o�o�o�o  DV�_z���� ���
��.�@�R� =v�a���������� �׏�*�mN�`�r� ��������̟ޟ�� ���8�J�5�n�Y��� }���ȯ�����A�"� 4�F�X�j�|������� Ŀֿ�ӯ���0�B� -�f�Qϊ�m����� ������,�>�P�b� t߆ߘߪ߼ߧ����� ���(�:�%�^�A�� ���ϸ������� �� $�6�H�Z�l�~���{� ������������ 2 Vh����� ���
.@R =O�s���� �/�*/</`/r/ �/�/�/�/�/�/�/?�?&?28�AGN_A�TC 1��K �AT&FV�0E02;AT�DP/6/9/2{/9p8ATA2>�,AT%G�1%B960k9�+++�?,�1H��?,�AIO_TY�PE  EC�/4?REFPOS�1 1� K x�O[H/O/ �O�MNO`O�O�O�O_ �OC_�Og__d_�_+K/2 1� KLON_��_o�_*o�_5A3 1��_�_�_ o�o�o|�o@oS4 1�Wo�io{o�o3W�oS5 1��o�oJ����jS6 1�����]�H���>�S7 1��(��:�t��ݏ���S8 1�����Ϗ	����r���)�SMASKw 1� O  
韜��ɗXNO�?���1.�8�1AMOTE�  �.DN�_CFG �U���5�0BPL_RANGQ��K!Y�POWER ��Q5 a�SM�_DRYPRG �%�%R���ȥT?ART ����UME_PROׯ��d�.D_EXEC_ENB  �5]�GSPD=�����Y3��TDB����R�Mÿ��MT_ѐT���S�D0OBOT�_NAME ��S�;9OB_O�RD_NUM ?���AH�80�0I$�	̗�s	�\������ ��e��	�@�}�D|��D0P�C_TIMEOU�T�� xD0S23�2n�1�Q; L�TEACH ?PENDAN��j��5��=Q�x0M�aintenance ConsK"�-��"+�t4KC�L/C�}�6���|� No Use�=[߹�F����NPO�ќ�5��_���CH_Lf@��U���	J�~�MAVAIL`����+��]�I�SPA�CE1 2�=L ����p���≢J@����8�?��� ���V� w�N������������� ���4�&G
l�} d	Q5U1��������� `4&G
l}Pd�#��2���� ����2A/b/@%/w/�//�/�3� ���	/�/-/O/^?�?B?�?�?�?�?�4 �/�/??&?�?J?l? {O�O_O�O�O�O�O�5�?OO1OCO�OgO �O�_�_|_�_�_�_o�6_*_<_N_`_o �_�_�o�o�o�o�o!�75oGoYoko}o +�o�o����)��>��8Rdv� �H�����ӏ%��F�-�[��G �N� R�;�
�� ����ԟ��� 
��.�@����c��� p���8�¯=�dؠ�� ϟ���!�3�E�W�i� _�q������x��կ ��'�9�K�]�oρ� w��ϛ���Ͽѿ��� �5�G�Y�k�}ߏߡ�����߻������ `S� @��8堯 F�"�*ل���� ��߇������,� ���V�h�2�<�N��� ����������.L 4v�R\n������
f�7�_MODE  ��^MS ���&����Ïb��*�	�&/�$CWOR�K_AD]	V���!R  ����t +/^ _INT�VAL]���hR_OPTION�&� h�$SC?AN_TIM\.��h�!R �(��30(�L8�"�����!��3��1�/@>.?�+��S22�41�9d�4�1"3��@���?�?�?���I-P���@����JO\OnOE@D� ��O�O�O�O�O�O_�_(_:_L_O���4X_�_�_��8�1>��;�o�� 1���pc]�t���Di�1��  � lS2��15 1 7oIo[omoo�o�o�o �o�o�o�o!3E Wi{����wc ���	��-�?�Q� c�u���������Ϗ� ���)�;�M�_�� �`[����ğ֟��� ��0�B�T�f�x��� ������ү�����$�7�  0��� o m��������ǿٿ� ���!�3�E�W�i�{� �ϟϱ�������v�� �/�A�S�e�w߉ߛ� �߿���������+� =�O�a�s������ ������ ��$�6�H� Z�l�~����������� ���� 2DVP�\�  �A���� ���%7I [m�����8��/ �/C (/N/`/r/�/�/�/�/ �/�/�/?F;/?�B?F�x1 �;?w=	1234�5678{�+�l�@�P�? �?�?�?�?O9/2O DOVOhOzO�O�O�O�O �O�O-/
__._@_R_ d_v_�_�_�_�_�_�O �_oo*o<oNo`oro �o�o�o�o�_�o�o &8J\n�� �o������"� 4�F�X�j�|������ ď֏�����0�B� T�f�����������ҟ �����,�>�m�b� t���������ί����(��6yI�[��@�`���������C�z  Bp*  � ���254F���$SCR_GRP� 1�(�e@(�l��0�@ `1 �[1s	 )�3�C� <�t�vrY�8P�}ϸkϤ����95C%����-u��ȡ����LR Ma�te 200iC� �190�1Շ0LR2C �3�=O���D�
f؜1u�2�U7��`1��v��@�u���	t����������$�^0� 2���_2T�gϡϊ�� o�F�D�f?��s������￶ht ,n�B�B˰�P�N�g�N�Aܰ�v�  @DЎ�N�@����  ?� ��J��H˰��y�N�F@ F�`������ A,Qwb�� �B��������B��_J� n�����/� %//I/��E+:3��6?|?�5��
�/�/�#��@=���?���6B�07�59�0@7���EL_D�EFAULT  �I����� ^1MIPOWERFL  V�xv5]2�0WFDOk6� v5 �ERVE�NT 1����O�t3C�L!D?UM_EIP?�8��j!AF_I�NEj0O�$!FIT�?=NOaO!Q�ΆO �PO�O!�RPC_MAINĮO�H��O�O�CVI�S�O�I��OE_!�TP8PPU<_�9d�4_�_!
PMON?_PROXY�_�6Ae�_�_XR�_�=f�_�)o!RDM_S�RV*o�9gouo!#RR8�o�4hdo�oK!
�@M�_�<i�o�!RLSYN�C4y8�oY!�ROS�?�|�4 H�tO�8c��� ��;��_�&���J� ��n������ȏڏ 7�I��m�4���X�����7ICE_KL �?%�; (%SVCPRG1�� ���!��3*�/�"�4R�W��5z��"�6�����7ʯϯ��C��5�9�� oG����o��� ���D����l��� ���񑼯7���_� �����4����]� ����������'�� տO����w��%ϟ� �M����u������ ����?�A��Ͽ�ђ �؟ꐊ���ɱ���� ����?�*�c�N��� �������������� );_J�n� �����% I4mX�|�� ���/�3//W/ i/T/�/x/�/�/�/�/��/�/?/??S?Ś_�DEV �9��MC:[8��im4OUT_R�f1~6i8REC 1q���f0�0 �1 	 �2�?�1�� �3OMO@O+OdO���
 �Z���6� s  UEBbf0K�q�0�0�f0Qʬ��2�3f0nf0��@ ��-�X�O�2Eb0��0'qE0_�O _�5"_�C&_L_:_p_ ^_�_�_�_�_�_�_�_ o o"oHo6oloNo`o �o�o�o�o�o�o  D2TVh�� ������
�@� .�P�v�X�������Џ �����*��N�<� r�`�������̟��ܟ ޟ�&��J�8�n��� b�����ȯ��دگ� "��3~A�(��P��� t�����ο�¿�� (��8�:�Lς�dϒ� �Ϧ����� ���$�6� �Z�H�~�lߎߴߢ� �ߺ������2� �V� D�z��n������� ��
���.�@�"�d�R� ��v����������� ��<*`N�� x����� 8HJ\������G�5V 1�&�< P_�1��AIO    i�0�=X>a?_TYP�E�?k2HELL_?CFG �z:f2�/ �B�/�/ %RSR�/�/�/ ?
?C?.?g?R?�?v? �?�?�?�?�?	O�?-O|?O/�  �!��@oO�O�O�C�I�A`PJ �N�A�@�W�gB2Pd�O�O�&H�K 1��+  �OE_@_R_d_�_�_�_ �_�_�_�_�_oo*o�<oeo`oro�oa&�#OMM ��/�o�"�FTOV_ENB�r$!}*OW_RE�G_UI�oe"IM/WAIT�b�I${�OUTv$&yT�IMu��`V�AL5's_UNI�T�c�v})MON_�ALIAS ?e~�i ( he! � ��$�6�Q&�c� u�����D���Ϗ�� ���)�;�M�_�q�� ������˟ݟ���� %�7��H�m������ N�ǯٯ������3� E�W�i�{�&�����ÿ տ習���/�A�� e�wωϛϭ�X����� ������=�O�a�s� ��0ߩ߻����ߊ��� �'�9�K���o��� ���b��������#� ��G�Y�k�}���:��� ��������1C U y����l ��	-�Qc u�2����� �/)/;/M/_/
/�/ �/�/�/�/v/�/?? %?7?�/[?m??�?<? �?�?�?�?�?�?!O3O EOWOiOO�O�O�O�O �O�O�O__/_�O@_ e_w_�_�_F_�_�_�_ �_o�_+o=oOoaoso o�o�o�o�o�o�o '9�o]o�� �P������s��$SMON_D�EFPRO ����:�� *SYS�TEM*  �l��*�RECAL�L ?}:� (� �}tpdi�sc 0=>la�ptop-u9n�qdgeh:59�28 cal_d�v.tp ove�r =>6320�94720:62?0723 5�͏�ߏ�s}tpconn 0 �������J�\��5cop�y virt:\�output\t�est.ls md:"�4�0���ӟ��}"ersrch� 0x160002��3 
���@�R� d�w�����-���Я���<z����� �� ������J�\��:z�f�rs:orderfil.dat	��tmpback\@���5�ƿؿ�1���b:*.*����8A ��=�O�a�t�xz�:\τ���0���,����}6z�a�ϔ� ���B�T���y���� /�����������ϭ� >�P�b�u���ϼ� �����τ��)߻�L� ^�q߃���9����� ����%��HZm� ����5������ �!��DVi�{��� 1��g��� �@/R/d/w
/� �/�/�/��/�/+<? N?`?s�/�;?�? �?�?�?'/�?JO\O o/�/?�/7O�O�O�/ �/�O#?�OF_X_k?}? O_3_�_�_�?�?�_ O�_BoTo�_yO_o �O�o�o�o�O�o�o-_ >Pbu_�_o�_� ���_o�)o�L� ^�qo�o9�ʏ܏ �o��%��H�Z�m ��5�Ɵ؟�� ��!���D�V�i�{�� ��1�¯ԯg������� /�@�R�d�w����-� ��п�������+�<��N�`�o��$SNP�X_ASG 1��������� P 0 �'%R[1]�@1.1f�l�?�o�%���Ͽ� ����� 6��@�l�Oߐ�s߅� �ߩ������� ��� V�9�`��o���� ���������@�#�5� v�Y������������� ��<`CU �y������ &	0\?�cu �����/�/ F/)/P/|/_/�/�/�/ �/�/�/?�/0??%? f?I?p?�??�?�?�? �?�? O,OOPO3OEO �OiO�O�O�O�O�O�O _�O _L_/_p_S_e_ �_�_�_�_�_ o�_�_ 6oo@oloOo�oso�o �o�o�o�o�o  V9`�o��� �����@�#�5� v�Y�������Џ��ŏ ���<��`�C�U� ��y���̟���ӟ� &�	�0�\�?���c�u� �������ϯ����F�)�P�|�_�x�PA�RAM ���}�� �	����P��p�OF�T_KB_CFG�  ����״PI�N_SIM  ��̶�/�A�ϰx��RVQSTP_DSB�̲}Ϻ����SR �	�� �& TEST �V����ԶTO�P_ON_ERR�  �����P_TN 	���A��RIN�G_PRM�� ���VDT_GRP� 1�����  	з��b�t߆ߘߪ� ���������+�(�:� L�^�p������� ���� ��$�6�H�Z� l�~������������� �� 2DV}z �������
 C@Rdv�� ����	///*/ </N/`/r/�/�/�/�/ �/�/�/??&?8?J? \?n?�?�?�?�?�?�? �?�?O"O4O[OXOjO |O�O�O�O�O�O�O�O !__0_B_T_f_x_�_ �_�_�_�_�_�_oo ,o>oPoboto�o�o�o �o�o�o�o(: Lsp�������� ��9�6�׳V�PRG_COUN�T�����d�ENB/�_�M��鴖�_UPD 1�	�8  
M����� ��-�(�:�L�u�p� ��������ʟܟ� � �$�M�H�Z�l����� ����ݯد���%� � 2�D�m�h�z������� ¿Կ����
��E�@� R�dύψϚϬ����� ������*�<�e�`� r߄߭ߨߺ��������\�YSDEBUG�n�Ӏ���d��"�S�P_PASSn��B?4�LOG ��΅�������
�  �����
MC:\`��a�_MPCf�΅����ҁ��� ҁ��S_AV �i���l������SV��TEM_TIMEw 1�΋ (u�Փq������T1?SVGUNSɀo��'�����ASK_OPTIONn��΅������BCCFG �΋O���I�2��`;A�I� r]o����� ��8J5nY �}�����/ �4//X/C/|/g/�/�/���,�/�/ ?? �/�/H?3?l?W?�?� �?��0�?�?�?O�? &OOJO8OZO\OnO�O �O�O�O�O�O_�O _ F_4_j_X_�_|_�_�_ �_�_�_o�X�  o2o Poboto�_�o�o�o�o �o�o�o:(^ L�p�����  ��$��H�6�X�~� l�����Ə���؏�� ���D�2�h�o���� ��ԟR�����.� �R�d�v�D������� ���Я����<�*� `�N���r�������޿ ̿��&��J�8�Z� \�nϤϒ���~����� �"�4߲�X�F�hߎ� |߲����ߤ������ �B�0�R�T�f��� �����������>� ,�b�P���t������� ������(��@R p������ �$6ZH~ l�������  //D/2/h/V/x/�/ �/�/�/�/�/
?�/? ?.?d?R?�?>�?�? �?�?�?r?OO(ONO <OrO�O�OdO�O�O�O �O_�O__&_\_J_ �_n_�_�_�_�_�_�_ �_"ooFo4ojoXozo |o�o�o�o�o�?  0BT�oxf�� �������>� ,�b�P�r�t������� ��Ώ��(��8�^� L���p�����ʟ��ڟ ܟ�$��H��o`�r� ������2�دƯ�����2��P��$TB�CSG_GRP �2����  �P� 
 ?�  {���w� ����տ��ѿ���/��A�T�[��b�d�0 �p�?P�	 wHBHA�L�͌�>@�B   C����0�ˀ��ϟ�D���ͣA���x���A��T8$�9��6ff��f�e@P�C�ώ�@�f����C��ߐ߮ߴ� ����%��%�D�W�"� 4���j�|�������?Y�����	�V3.00s�	�lr2c��	�*2�*�O�A� ��ѳ�33P�d��� 8x�J�y�  �������T�JCFG -��l� o���+��������=K
%�K q\������ ��7"[F j������� !//E/0/i/T/f/�/ �/�/�/�/�/s���? ?(?�/[?F?k?�?|? �?�?�?�?�?O!O3O �?WOBO{OfO�O�OP� <��O��O�O�O0__ T_B_x_f_�_�_�_�_ �_�_�_oo>o,oNo Pobo�o�o�o�o�o�o �o:(^L� �����h� �� $��H�6�l�Z�|��� ��Ə��֏؏� �� D�V�h�z�4����� ��ҟԟ��
�@�.� d�R���v�������� Я���*��:�<�N� ��r�����̿���޿  �&��>�P�b�ϒ� �ϢϤ϶�������� 4�F�X�j�(ߎ�|߲� ������������B� 0�f�T��x���� �������,��P�>� t�b������������� ��&(:p^ ����t���� �6$ZH~l� ������/2/  /V/D/z/�/�/�/j/ �/�/�/�/?.??R? @?v?d?�?�?�?�?�? �?�?OO<O*O`ONO pO�O�O�O�O�O�O_ �O__&_\_�t_�_ �_B_�_�_�_�_�_"o oFo4ojo|o�o�o^o �o�o�o�o�o0B �oxf���� �����>�,�b� P���t���������Ώ ��(��L�:�\��� p�����ʟ��� ��_ �*��_�l�Z���~� ����į�د� �2� ��h�V���z���¿ Կ濠�
�����.� d�Rψ�vϬϚ��Ͼ� �����*��N�<�r� `߂߄ߖ��ߺ����� ��8�&�H�n�\�� �>�����x������ 4�"�X�F�|�j����� ����������
 Tfx�D��� ���P> tb������ �//:/(/^/L/n/ p/�/�/�/�/�/ ?�/ $?6?��N?`?r??�? �?�?�?�?�?�? OO DOVOhOzO8O�O�O�O8�O�O�N  PS� V$_R�$�TBJOP_GR�P 2��E��  ?�hW<RCS�J\��@O0WP�R@T^�P � ��T�T� �Q[R	 ��BL  �UCр� D*W[Q�_�_?�fffe:l�B �P�ff@�`�33D   $a�U3o>g�_�_po�l��P�e9<�bbY��?٪``$o�o�UA��gD�`$��co�Quz9��P�Aa�P@a���C�Z`Ep�o]�A6ffpu`aD/�U�h�͔r��~ �a�RieAq�`�q��!@9q�|�d&`%����c333D�\P8o���?�`?L�pAp[QB�b�k�}� ���z�� >�ffԁL���T�f�� fo ��Nw@�*�8�f� ��r�,���П��ȟ�� '����F�`�J�X���,��SC�Vء��	V3.00�S�lr2c�T*���TQ�� �E���E�A �E��E��3�E�iNE�!h�E�فEۑ��E�I�E���E���E�r�F�F��FM(F�5�FBFaO�F�\F"f�,�z  E�@ �E�� E�� �E�  E������ E����� �EȆ�Ԏ�ᆰ��� F   F�� F$ Fj�` F�@ F��P F�` 9��IR9�o��D�L�_ ��V���LQ�8TESTPARS�XUP�9SHRk�ABLE� 1�J[4�SDV�+� �0�V�VȡV�WQV�	V�
�V�Vȥ�QV��V�V�뱅�RDI��TQ�϶���������f�On߀ۊߜ߮�H���ކ�Sl�RS 0� ������������� #�5�G�Y�k�}����� ��������/]k�o�� *	�%�7�I������+�=�O؆�NUM�  �ETQ��PP �밆�_?CFG �����Q@<PIMEBF_TTq��RS~�;GVER�<Q;�R 1�J[
 8I�RP� �@5  ����� �//&/8/J/\/n/ �/�/�/�/�/�/#?�/ ?Y?4?F?\?j?|?{�_�h@R
<PM�I_CHANG �R �3DBGLV�Q`IR;Q�0ET�HERAD ?*�E;@�S �?�?xTO6V�0ROUTe!JZ!�D�OwL?SNMASK0HRS>AA255.�E���O�O8TOOLOF/S_DIq��5I�ORQCTRL C�s[���n]8]_ �_�_�_�_�_�_�_o "o4oFo�
�_Tofo�o�g�PE_DETA�IH3ZPON_S�VOFF)_�cP_?MON �"P�2�iSTRTCH/K �J^mO�b�VTCOMPAT��h;C�d�`FPROoG %JZ%j��=?qqISPLA�Yr��j_INST+_M�@ �|�g�t�USe]orLCK���{QUICKM�E�0)�orSCRE�F�3Jtps��or�a�f��2w��_{���ZyISR_�GRP 1�JY/ ؛ 6� ����;�)�_�M��8����Y������ �͕�����/��S� A�w�e�������ѯ�� �����=�+�M�s��	123456�78����f�X`�1��Ћ
 �}i�pnl/۰gen.htm������0�B�X�Pan�el setupF�}<�ϘϪϼ����� u�k��*�<� N�`�r��ϖ�ߺ��� ������ߝ�J�\� n�����I�?��� ���"�4�F���j��� ������������_�q� 0BTfx�� ����� >�bt����|3�~UALRM�p�G ?J[
  �*/!/R/E/v/ i/�/�/�/�/�/�/�/�??<?�SEV � �n6�E?CFG ��m�6���A�1   B��t
 =?�s3E�? �?�?OO+O=OOOaO�sO�O�Gz1ʂ��k� SΟ�OH7Isv?}{�`(%0?"_p_ I_4_m_X_�_|_�_�_ �_�_�_o�_3o�L�c �M�OAoI_E��HI�p1��i  �( k`���(/SOFTPA�RT/GENLI�NK?curre�nt=menup�age,153,�1}o�o&�'�o�n3�op���5G�b71`����+��q+��eed�it�bCAL_DAV�}�����0�)C�U�TESTl�����#�5� �o�,148,27����������)oߟ���'�9� ȟ]�o���������è�R��aR����%� 7�I�L�m�������� ǿV�����!�3�E� Կ�{ύϟϱ����� d�����/�A�S��� w߉ߛ߭߿���`�r� ��+�=�O�a��߅� ��������ʯܯ� '�9�K�]�o�r���� ��������|�#5 GYk}��� ����1CU gy����� �	/�-/?/Q/c/u/ �//�/�/�/�/�/? ���;?M?_?q?�?�? �/�?�?�?�?OO�? 7OIO[OmOO�O�O2O �O�O�O�O_!_�OE_ W_i_{_�_�_._�_�_ �_�_oo/o�_Soeo wo�o�o�o<o�o�o�o +?(?as� ����o���� '�9���o������� ��ɏX�����#�5� G�֏k�}�������ş T�f�����1�C�U� �y���������ӯb����	��-�?�Q�<���$UI_PAN�EDATA 1��������  	�} � frh/cgt�p/wholed?ev.stmc����ӿ����)  ri��.�Ip��F�X�j� |ώϠ�ϲ��Ͻ��� ���0��T�;�xߊ� q߮ߕ��������Bv���  �  
is$ @�E�W�i�{����� ��6�������/�A� ��e�w�^��������� ������+O6 s�l�� ��� ������1C �g������ �L	///?/&/c/ u/\/�/�/�/�/�/�/ �/?�/;?M?���? �?�?�?�?�?0?Ot %O7OIO[OmOO�O�? �O�O�O�O�O_�O3_ _W_i_P_�_t_�_�_ �_�_Z?l?o/oAoSo eowo�_�o�o O�o�o �o+�oO6s �l������ �'�9� �]�D����_ o�oɏۏ����#� v�G��ok�}������� ş,�������C� U�<�y�`�������ӯ ����ޯ�-�����c� u�����������T� ��)�;�M�_�q�ؿ ��|ϹϠ�������� ��7�I�0�m�Tߑߣ� ����:�L����!�3� E�W��{�� ϱ��� �������r�/��S� e�L���p��������� �� =$a����}�r�����)�*��V hz����� ���.//R/9/v/ �/o/�/�/�/�/�/?��������$UI_�PANELINK� 1����  �  ���}1234567890_?q?�? �?�?�?�4��]?�?�? OO1OCO�?gOyO�O �O�O�OYIY0:�M���[0  SOF�TPART/GE�NA1?CONFI�G=SINGLE�&PRIM=mainedit �O�I_[_m_YJ_$_M=�wintpe,1 @_�_�_�_�]�_$o6o HoZolooo�o�o�o �o�o�o�o
2DV hz����� ���.�@�R�d�v� �� �����Џ���~�M 0,  9P E=Por?S�5�co:�{�^������� ͟ߟ��'�9�� ]�o�R����O�O���� �Z1�/�%�7�I�[� m�`C�������Ϳ߿ 񿀿�'�9�K�]�o� �L���э͙�S���� �������#ߒS;�M� _�q߃ߕߧ�6����� ����%��I�[�m� ���2��������� �!�3���W�i�{��� ����@������� /��Sew��� �.���|�# G*k}`��� ���/�1/C/֤ �͡�ۯ}����/�/�/ �/�/?�2?D?V?h? z?�??�?�?�?�?�? 
OO�ϝϯ�dOvO�O �O�O�OE�O�O__ *_<_N_�Or_�_�_�_ �_�_[_�_oo&o8o Jo�_no�o�o�o�o�o �oio�o"4FX �o|�����e ���0�B�T�f�� ��/���������ُ ���>�P�3�t���i� ����Ο��O/�s/(� �/L�^�p��������� �?ܯ� ��$�6�ů Z�l�~�������#O5O GO�� �2�D�V�h� ��Ϟϰ�������u� 
��.�@�R�d�v�� �߬߾������߃�� *�<�N�`�r���� �����������&�8� J�\�n���������� ������m�"4ßX jM�q���� ��BT7x ������A��/ /,/>/P/C�t/�/�/ �/�/�/�/o/??(? :?L?^?Ϳ߿�?�? �?�?�? OO�?6OHO ZOlO~O�OO�O�O�O �O�O_�O2_D_V_h_ z_�_�_-_�_�_�_�_ 
oo�_@oRodovo�o �o)o�o�o�o�o *�oN`r��� ��m��&�8� �\�n�Q���u���ȏ ������"���?�?��{��$UI_P�OSTYPE  ��5� �	k�{��_QU�ICKMEN  ���j�����RESTORE 1ו5�  ���/
�2�D�h�m c�������¯ԯw��� 
��.�@��d�v��� ����W���˿ݿO�� *�<�N�`�τϖϨ� �����ρ���&�8� J���W�i�{��϶��� �����ߡ�"�4�F�X� j���������� �����y�+�T�f�x� ����?��������� ��,>Pbt�� ����( �L^p���I���� //��SC�REܐ?��u1sc-�uU2M$3M$4M$5M$�6M$7M$8M!��UGSER/ 4/F"T. �O#ksW#�$4�$5*�$6�$7�$8�!���NDO_CFG �؜�  ,� ���PDATE ��)�Non�e V��SEUFRAME  
���&,1RTOL_�ABRT7?��N3E�NBX?I8GRP �1�!��Cz  A��3�1��?�?�?�?�?FO"OG:�ېUx81g;MSKG  {5�Ag;N41%a��B%��O���VISCAND_wMAXyEI�c8��@FAIL_IM)Gy@f���#�8�@�IMREGNUMryG
�KRSIZyC�,���$,SO�NTMOUW0{D��%�VU�#�c�� �P�2F�R:\�O � �MC:\XS\wLOG�VB@4 !�O�_�Q�_o
��z MCV��_�SUD10fE�X9k
�f�wV�2�ꜙ�p(��=��͓o��j�o�o�o �o�o�o�o 2D�Vhz��KPO6�4_?S�0��n6�uQ0LI Q�z�xr�qV� �|f@�w��� =	�xSZ�V�~����wWA�I��DSTAT ܛ;�@�_ď֏��$����EP12D�WP  ��P G/����q�AP-���B_JMPERRw 1ݜ�
  � �2345678901�������ʟ�� ϟ��$��H�;�l��_�q����LT@MLO�W���P�@�P_TI�_X�('�@MPH?ASE  53���CSHIFT�UB1~k
 < ���Ob��A�g���w� ��ֿ��������� T�+�=ϊ�a�s��ϗ� ���������>��'��t�K�!��#ޛ:	�VSFT1�sV:�@M�� �5��4� �0��UA�  �B8���Ќ�0p������Ҫ��e@��ME*�{D�'���q��W&%�!�M�$�~k���9@�$~�TDINENDcXdHz�AOx@[O��aZ��S�︕��yE����G ����2�������<���RELE�y?�w�^_pVz�_ACT�IV���H��0A ���K��B#&��R�D�p��
1YBOX� ��-�����2�D�1�90.0.� 83v��254��2�p�&���robo�t�ԟ   �pN g�pc� �{�v�xx���$%ZABC�3�=,{�낆;- !/^/E/W/i/{/�/�/ �/�/�/?�/6??/?$l?!ZAT����