��   �A��*SYST�EM*��V7.7�077 2/6�/2013 A� ���$$CL�ASS  �S��(��D��D VIRTUAL%�7MNUFRAM�E AF�D� � 	� 88�?� ��}��y���� ��1=gQ s������	/��/?/��WNUM  ��>l�  �WTOOLa4 
wY/�/5/�/�/ �/?5??A?k?U?���t5s?  Bo��^�1C  G __? �?�?]?�?OO%OOO 9O[O�OoO�O�Og,�!
{&���'* 