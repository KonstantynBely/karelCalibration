��   ��A��*SYST�EM*��V7.7�077 2/6�/2013 A�   ����DRYRUN_T�   � $�'ENB  �$NUM_POR�TA ESU@�$STATE �P TCOL_��P�MPMCmGRP__MASKZE� �OTIONNLO?G_INFONi�AVcFLTR_�EMPTYd $PROD__ L ��ESTOP_DS�BLAPOW_R�ECOVAOPR��&J_  �4 $TYPE�NFST_IDX؞$_ICI � �MIX_BG�-� G_NA�Mc %$MOD�c_USdkIFoY_TId K�MKR-  �$LINc  { �_SIZ��K� ?.  �$USE_FL�GA���i�S�IMA�Q�QB�
'SCANzAX�'+IN'*I��_C7OUNrRO���3!_TMR_VA�g�h>� i��'` ��&pܸ!�+WAR�*��$$CLAS�S  �����!��5��5� VIRTUz �/� '/ �
55���*����C80�!�J5��5I1&; ��?�?�?�?�?�?�? O!O3OEOWOiO{O�O`�O�Oc?+ W?
5{01 ��X�O__  W1J0��C O 1&;G 4%�On_��G1 W1\_�_�_�_�_�_�_ o�_1oCo"ogoFoXo �o|o�o�o�oW1@S��&=^9J0�� -rJ16t,G1
1>q�o `r������ ���&�8�??�c>q W1j�|�������ď֏ �����0�B�T��$�?T�1&9 K������ӟ� ��	��-�?�Q�c�u� J�������̯ޯ�� �&�8�J�\�n����� ����ȿڿ����"� 4�F�X�j�|ώϙ��� ����������0�B� T�f�xߊߕϧ����� ������,�>�P�b� t���߼������� ��(�:�L�^�p��� ������������  $6HZl~�� ������� 2 DVhz���&V