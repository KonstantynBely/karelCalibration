��   &��A��*SYST�EM*��V7.7�0107 10�/3/2018 A   ����DMR_GR�P_T  �� $MA��R_�DONE  �$OT_MINUS   	G�PLN8COUN:P T REF>wKPOOtlTp�BCKLSH_S�IGoSEACH�MST>pSPC��
�MOVB RA�DAPT_INE�RP �FRIC��
COL_P M�
GRAV��� �HIS��DSP�?�HIFT_E�RRO�  �N\ApMCHY Sw�ARM_PARA�# d7ANG�C M2pCLD�E�CALIB�� DB$GEA�R�2� RING���< �PLC�L* ��ST�A� mTRQ_M<��LINK"2&�SX<*Y<*Z/)I�I*IW*Ie$ �R�V* L $� ENBpV_D�EBU��!PN�U;%� UNEVE�ox�!8� �$��ASS  �����!������ VIRTUAL��/1' 1 5�� 
��� ��b?M?�? q?�?�?�?�?�?O�6�H+O�71HO6M,�����w����R�.A��E?�# (.�5O�O 1O[L�O�O�O�O�O_�KA_GR0_m__j_�_��d�_�_�_�_���=L���_"o?�#o��@�Cohozo�o �o�o�o�o�o�o
.�_ 5YgwQ�4  2�_�� �� ��$�6�H�Z���<���������̏ ޏ����&�8�J�����$% 15B1D�U5a�� ���_���_�ϟ�� ,��)�b�M���q��� ����ݯ�����(�� L�7�p�[�m�����ʿ ���տ߯!��H�߿ l�Wϐ�{ϴϟϱ��� �����2��#�e�'� ��#߰ߛ��߿����� ��.��R�=�v�]�g� ��k���g������� <�'�9�r�]������� ����������8# \G�k}��� �����1�X� |g������ �/	/B/)/3u/7/ �/3/�/�/�/�/?�/�?>?)?b?M?�?[�R5Vk�r�`{?�?s?�?Hjx�?&O8OJO \OnO�O�O�O�O�O�O �O�O_"_4_F_X_j_ |_�_�_�_�_�_�?�_ o�_0ooToOxo�o �o�o�o�o�o�o ,>Pbt��� ������(�:� Ao^�I�n���{���ko ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯�����߯ �Ϗ@�R�d�v����� ����п�����*� <�N�`�rτϖϨϺ� �������	�&��J� 1�Z߀�3��߶����� �����"�4�F�X�j� |������������ ��0�B�T�[ߕߊ� u����������� ,>Pbt��� ����(: L^p������ ���/�6/��Z/ l/~/�/�/�/�/�/�/ �/? ?2?D?V?h?z? �?�?�?�?�?�?�?
O O#/@O+OdOvO]O�O M/�O�O�O�O__*_ <_N_`_r_�_�_�_�_ �_�_�_oo&o8oJo \ono�o�O�o�e