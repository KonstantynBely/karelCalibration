��  ë�A��*SYST�EM*��V7.7�077 2/6�/2013 A�Q  �����ABSPOS_G�RP_T   � $PARA�M  �  �ALRM_�RECOV1   $ALMO�ENB��]ON�iI M_IF1� D $ENA�BLE k LA�ST_^  d�U�K}MAX�� $LDEBU�G@  
FPC�OUPLED1� $[PP_PROCES0 � ��1����URE�Q1 � $�SOFT; T_I�D�TOTAL_�EQ� $,N�O/PS_SPI�_INDE��$�DX�SCREE�N_NAME {�SIGNj���&PK_F�I� 	$TH{KY�PANE7�  	$DUM�MY12� �3��4�GRG_S�TR1 � �$TIT�$I��1&�$�$T�$5&6&7&8&9'0''��%!'�%5'1?'1*I'1S'1]'2h"GSBN_CFG1 � 8 $CNV_JNT_* ��DATA_CM�NT�!$FLA�GSL*CHEC�K��AT_CE�LLSETUP � P� HOM�E_IO� %�:3MACROF2R�EPRO8�DRUeNCD�i2SMp5�F�AUTOBA�CKU0 � }�	DEVIC#sTIh�$DFMD�ST�0B 3�$INTERVA�L�DISP_U�NIT��0_DO��6ERR�9FR_�Fa�INGRkES�!Y0Q_�3t4C_WA�4�12H�GX_D�#	 �d $CARD�_EXIST��$FSSB_TY�Pi� CHKBD�_SE�5AGN G�� $SLO�T_NUMZ�AP'REV��G �1�_EDIT1
 W� h1G=H0yS?@f%$EP�Y$OPc ��0LETE_OK�zBUS�P_CR�yA$�4�FAZ0LACIwY1KR�@�k �1COMMENy@$DGV]QP�� ���AL*O�U�B , $��1V1AB0~ O�L�UR"2CAM_�;1 x�f$ATTR��@0�ANN�@�IMG?_HEIGHyAc�WIDTH�VT�CYU�0F_ASwPECyA$M@7EXP;$� Mf��CFcD X O$GR� � S!1zU`BfPNFLIC`<~d
UIREs3���AOMqWITC)H}cX`N.0S_d�S�G0 � 
$WARNM'@f�̍@� LI? �aNS=T� CORN��1�FLTR�eTRA�T@0T�`  $ACC�1"p '|�'rORIkP�C�k;RTq0_SF� �!�CHGI1 E[ Tz`u3IPpCTYVD�@*2 �P��`� 1zB*HD��SJ* ��q2�v3��v4�v5�v6�v7��v8�v9�vqO�$ <� so�o�h��s1�PO_MOR~. t 0�Ev�NG�8`TBA� 5c���A�����]@����ϋaP�0Ѕ*��h�`
P�@�2� �,p�J,p_Rrrqo@+�1J/r/�J�JVq@��Cj��m�g��ustP�_}0OF� 2  @� RO_���Wa�IT8C��NOM_�0�1ەq34 ��cD� �;����hP���mEXpG�0� �F�p%r
$TF�x�JF�D3ԐTO��3&@U=0�� e�H�24�T1��	E�� �e��f�t�f���DBG;a�� k@$�PPU8�3�f):��&A�AX 1�dUN�$;AI�3BUFuF����! |�`��`[PI��Pr�EMq�M~�䠁�Fr�SIMQS��G�`�QE���F��MC{�k �$}1JB�`S�}1DEC���������x� ě0CH�NS_EMP�r#$Gg�=Ǎ@_��q3�
p1_FP󔞡TCh�@`�b��q0�c}�y�G�� V�AԂ�!!���JR!0ԂSEGGFRA.pv 7aR��T_LIN�C��PCVF������Y ���Q��)B����( '���f�e �S���Q��.0�p�B�8�A����SIZC����z�T��g������QRSINF3��p�� ��?�������؉����Lot��G�*�CRC�eFCCC�`+���T� h��mh�SbA��h�*��f��:�D�d�c��C��PTA����w@��L����EV���jF��_��F��N&�G�� �X������1i��! ��,��h#RGNP��0qF���R�}�D���2}�LEW N��Hc6���C�K�۲}RcDx :�@L��ou2���A6N`�Co�$LGp��B@�1aP��s@�dWaA?@����~0R���dM�E%`��d�_RAs3dAZC���z��OkqFC�RH`X`F�`��}��,�ADI ;� 6b� ���` �p�`5cn�S�@1�L7a�AMP���PY8C�U�MwpU��iQU� $�P��C�C�G1������DBP�XWO����p�$SK��2!�DB]T TRL�1 ���Q0Ti� �P�DJ��4LAY_CAL`�1R !'PL	3&@�0ED�Q5'�Q5'"̡���1!�W�;PR� 
�1� 0�1" �PA�$�q$�� ��L�)#�/�#mp�0$��/�$C�!%�/�$E3NEqr�&�/�#�d REp�"'H� �O)@"$LF3#$�#xB� W;4���FO[ _D0m�RO(@���u��j��~�3RIGGER�6�PA%S���ETUsRN�2RcMR_���TU�`?�u0EW5M����GN�P���zBLA��E��$�$P#�CP� ��&�@�Qk�C5D�mpD��A#�p4\1i�FGO�_AWAY�2MO���fQg�CS_n(<�QIS  ����c�C���A����B�t�Cn��A"r�FW���DNTV@��BVkQ�����S˳W��sU�J&�U�� ��S�AFE�ZV_SV>6bEXCLUl������ONLA��SY���Q�tOTBa��H�I_V/M�PPL�Y_�a��VRFY�_#�q�Bd�_ #)0���_+�Ipg `"�@SG3� *�b݀�0 AM�@��a*����0��Vi|.b%fANNUN� ,rLdIDp�U�2~S@�`mijarj�f���堫@I�"+��c$FOb�׀OT@�w1 $DUM�MY���d[!�d١��& �E, ` 8�HExs��b�S|B$�SUFFI��@ ��@�a5��g6�a(�DMSW�E- 8��KEYI����TMZ1^ӌqL�1�vIN������. D��HOST? !�r���t�[ �t٠�tYp�pEMp>���$��SBL��;UL��/ �|�3����T50�!0 ϴ $9��ESAMP�ԕF���������I�0��$SUBe�Q�� �C�:��G�SAV��r����G�C� ˇ�PnfP$�80E��YN_Bn�1 0��DIadb�@O���}$]��R_I�� �E�NC2_ST � 2
ԇ J���L�q~S# :����!3�M��I��1:�p�4 � L�3�M��0�0K�4'a��AVERp�q��}�M�DSP�v��PC�U����\ì�VALUŗHiE� ��M�IP@����OPP7  �T!HS ���6�S�F�F􁳠dL�0�T���SC�Q�d:�E�To�5zrFULL_DUY�da�0��0O�w�h�OT��~�0NOAUTO�!6�p$�\���c�l�
�C` �CL���z���L�� 7H *�AL���n�b���$�0 P�˴��ֲ��[!���a���Yq��dq��7��8J��9��0����1��U1��1��1Ⱥ1պU1�1�1��2
ʩ2����2��2��2�Ⱥ2պ2�2�2*��3
�3��3����U3��3Ⱥ3պ3�3�3��4
�iq��;SE�"8 <��~��`�;I�����/���QFE�0�0� 9 �,��Q?hpz@^ ?Q�А��ER@B#� ��@��� :�`�$TP�$V�ARI�<��UP�2�P; �pq�TD ��S|�1`3���iq�r�BAC�< T�pr��)��bP�P o�IFI)�P ���TU���P���F�0|��� =t ;'�0Ԡ��P'�ST(&�� HR&�r0E����	
%�C��	���_Cr��N�r��B��p�h�FO�RCEUP%bn�FWLUS�`HN �xE�h�RD_CMK@qE(����IN_��&vPg�REMM�F ~Q��M �� 3
�K	N0�EFF���N@IN�A��O�VMl	OVAl	TgROV���DT��mDTMX���m {@�
��? �*[ ��CL��_:p']@d$�-	_
�;_T��TX
��@AQD� ��}��}!V1�� RQ��LIMI#T_�a椀�M��sCLmd}�RIV	��a��EAR��IOF*PCC�����B�B�g�CM@��R ��GCLF�G!DaYM(/�aR#5TWCDG��| s% �sSS& �s> P�a(�!r1��wP_�!�(J�!1��E�3�!3�+=5�&�GRA����?w��kPW��OyNT��EBUG)S�&2*�P{@a�_E �@�P�Q�S_�TERMB5AK5���ORI�G0BK5�O�S#M_�Pr�G0CK5~@��TA�9DK5���UPB�E� -�zAa�@.PY3.@A�$SEG�:f EL�EUUSE�@NFI,��2�1ޠp4�4�B$UF6P�!$�FQ4@�wAG�0TQ�&�HSNST� PATm�piBP'THJ�AߠE�p� �2�P؀	E)�؁��1�R�@�InaSHFT�_��1oA�H_SHOQR ܣ�6 �0$�7r�@Dq�'�OVR#��na�@I�@�U�b �QAYLO=�z���I'"�oAj�!�j�ERV��:Qh��J��OG� @�B0����U>���Rz!P"�ASYM.��"��1WJG�уE S�A�YvR�U�T @ ���E)�ᥳEP!�WP,!�WOR @MB��_GRSMT�F�cGR��3laPA.@���`�q�uG � u����TOC�1��`P�@ �$OP@��ဝpՓá ��YO��RE�`RCb�AO�pтpBe�`�RmE u�h�A��e$7PWR�IM�ekR�R_�c4��qB �H2H���p_AD�DR��H_LENAGqByqnq�q�R��]S�I H��S�� �q0Ӧu>Ӵu���u��#SE�'�LrS��J $N�`��_�OFF��rPRM�� �HT�TP_�H�K (^pOBJ?"ip��[$��LE`C!�>ȠL � �׬��AB_~TS�s�S�{`��*�LVN�KR���eHIT��BG��LO�qt�fN�`͂���`���`SS{ F��HW��A�M�p}`INCPU�"VIS�0�����+��t,��t,��� �IWOLN��N̠��C��$SLQb���PUT_�$��`{�P �V���F�_AS�"O��$AL��I����A��U�0��@�af��`q�<PH�Y���Ó![���U9O��#P `�������ڔ� �2�pP ���`(�L��Y�B�D���UJ�Q�z�N�EWJOG-G��DISx�[�K-�f�#�R 
�WAV�ǢC�TR�CǢFLAG��"[�LG�dS �����Y�3LG_SIZo���������FD)�I�4�E� *��D0���c$��� 𖶦���K���D0��� SCH_��߅p��2��N��F�T����E�"~�������U�
�
�{`L�	�DAU/�EA�-��dE��;�GH�bt���BO}O��Uh Aɒ���IT��y�[0ŖR;EC��SCR�𙃖ʑDIēS.@��RGO���˒����d��$����SU���W�Ĳ��Ľ�JGM$�MN�CH,�FNKEuY%�KM�PRGK��UFY�PY�FWDvY�HL��STPY��VY�@Y؀�Y�RS"��H1`uۺ�CT�� �R��� �$�U	�m�@��
R�ݠғ`�G=ن�@POd�ڻŦ�M��FOCUd�RG�EX��TUIK�I{�����	������I�M��@A�S�`��p�@������ANA����2�VAILl�C�L!�UDCS_H!I+4`�s_�Oe�
!"h�S���|�S����IGN4��F�J��9T�be�_BUj � �V !PT�$�*��rv�Ϥd�@�A
VrW !Pi�'��T�0�1?2?3?�_� X � �i�=a�5���Ņ�ID$� tbP5R�bOh �Ĭ\A�ST	�RF�Y�� �@�  W$E�C�y�����FFLa�� Y L�؟0��@���`�qFtǀ�FwҬ�_ Z i`�����b���>0C��[ =�p CLDP	��UTRQLI{��T����FLG�� 1��O�D�����LD8���ORG���� ��hW>(�siT�r� 4\ �#0��վJ�Sy`T�70#0�' �$�!�#RCLMC�$B/T/�)Q��!=19I�p_d] d��RQ73$DSTB��p�   6��-8A�X�R /8I<EXWCES�bz 5Mp
�1^��2�T�2���0_�p"6_A@:&��;G?Y80K�d�` \�GROU���t$MB �LI�9�CREQUIR�DB�aLO#KDEB�Ur� 1LYM��a@gbʑ`@�C�" 1#ND��`c`b����̨�CDC���IN�'��C��Z`���H��N���a#�� �EPS�T�� c\rLOC�RITp��P��Ap�1 1ODA�Q��d X��ON�cF�R�fV�	Xಐb�U���w �F�X0IGG�� e �y X�a��X4�XR�Q%��Y�	��X	��V�0ғDATA$`E�a��a��N��f t W$MDEaI:�)Sf��^d�![gH5P�@]exz��a_cANSW�aP^d�a��^eD�)AR�z�� Xpg �0C�U4�V�`�=URR2{�h D2�`A���A�! d$CA�LI&0��GS�w2NK�RINb�t<�'NTEg�(i�bCu���=RBqg�_N�qj@Pukr���$ht�2kuy7DIV�&DHi0jp:+�l $Vp�Cv�$M�$Z0R�<!T 0R���b�em�H �$BEL�T˪ZACCEL���;�"�IRC�O�݁m��T����$PSi0�Lt� ڰW��Cp8��T�9�PATH���.���3]��Pl1_<�r���Ł�"S Cr��_M=G��$DD�9���$FW�`7`����.���DE�P�PABNe�ROTSPEEՂ@L� �JN�@��(0�t��$USE_p�P�&�ܦSY>��p�! ��QYN0A����OsFFua��MOU߁3NGJ�܀OL~�ٔINC�d2Q��-2x��� -2ENCSp�a2U��+4R�IN��I]�B����"n�V�E��s^�23_UyPօp�LOWL��A[�` '���D>�@2@Ep]'��2C[p�W�MOS���4MO���0�'PERCH  ��OV����� �������$�8S+� � 2@������V�0^�O�L�P��7O�U��UP"�������TR�K��AYLOA �J��1��]�͵³3P� �RTI�1	�� MO�O�-2�28 �`4�wٳ��?�p�DUM2��S_BCKLSH_C]� P�ϐΦ����bn�"��y�Ñ���CLAL� V��!��� ��CH�K �SՐRTY@����C�
*!6a_�Nä_UM����C����SCL�W�LM?T_J1_L< 0-օa:�E4�U�G�pD�J�P�J�SPCd�0ȑZ���3�PC �3�!H_A@���C� csXT���CN_rN���.�S��%�V���:����]�9�2��C' �SH�r �*�*!9�9� p��^����9���PA���_	P��_�"�Ŷ�0!ճ����JG�����~�OG��,�TORQU��ON��޹*�`B٢-�*�L�_W���_�sj��sj��sj�UIr�I��I�sFKP�]�J�!��c!�VC"�0'4�2��1��{08��82��JRK��+�� DBL_SMt���"M�@_DL�q�"GRVq�j�sj�sKH_��I���
�COS��LN - �����p�	�p�	 �����FZ� ٦�KMY�D�TH|�eTHET0��NK23�s��s� [CB�CB�sC&1�n2�����s��SqB�s��GTS�1W�C.�2Q�����$x�'3$DU�� �8A!r��2P&��19Qb8V$NE�4�PAI� ���"%�v$�p�A��%�'����LPH�5�"h��"S ��3�33�"+3(:2�pV�(V�(�p��,V�*V;V;V�";V0;V>;VL9H��(�&�2�-n�H;H�;H";H0;H>;H*L9O�,O�(O}I�.UO�*O;O;O";UO0;O>;O2F�"�Y�T�'SPBALANCE_T�@SLE�H_�S�PHq�hR�hR3PFULClX�R{W�R�3Uz1i
�UTOy_����T1T2�Y�2N���`��Tq@���Ps d���T��O�p!�L�INSE9G���REVf���Q�DIF��zy1jl_g�r1k��OBUa��t$yMI`���S?LCHWAR>���AB��u$ME�CH�Tˑ�a��AX˱Py��f�'�r�P�l 
�bI��:�ROB�CRW�-u��=(�pMSK_KP�t_n P �P_��AR��r_tn���18�c�a�_p`�y�_p�aI�N:a�MTCO�M_C���po � ݀g`4�$N'ORES��r��`�rop 8U�GRJ��eSD� ABג$XYZ_DA�!<F�r�DEBU:a�q����pq _P$��C;OD�� 1�����`��$BUF/INDXa�Hp"��MORRsr $�qU&���u��ӑyçDB:!��bGi�s� � $SIMUL��8��>���F��OBJEjP��AD�JUSψAY_	I��8�D���s�Ԑ�_FIב=s�T Z��c����`b�"��(�b`p0G�D��FRiIW�d�Tg�RO%��A�Eb�
HpOPsWO> Vpt0>��SYSBU0[�$�SOP��I�����U<��b`PRUN�rڕPArpDٖ�b��1�_OUTΑ�a�t{$�IMAG��i\pv PDaIM���1�IN[ �0�RGOVRDY�˒���aP�/�a�� L_�P0B�}����RB�� e��MkᜪEDb�*�` �N�@M��~�o)*�\�SLjP�Vpu x $OwVSLfSDI��DEX���q�����$o��Vb��N�A�@�'��,�'�D�M~�z��]�_SETK�Vpv @U�^��e�p�RI��j�
q�_�}�����Hpdà>*� w H\q�`���ATUS<�$�TRCx T�X�ѳBSTMڷıI��P��4}Ѱ���Vpx DB\pE���β�0Ehb�ϱ�����ϱEXE�հ����)�=��f�y�m�]p԰UP�L�9$�`6�XNN����x������ �PG�u7zWUBñ�e���ñ��JMPWAeI[�P���LO7��FA`��$RCVFAIL_Cwq����R9��p�c��(��}�"�-�AR_PL��DBTB��,⾐gBWD ��pUM*��"�IG�7��Qc�T#NLW�"�}�Ry�iӂ��E�����Hp��D�EFSP` {# L\p�`��_��Ճ��UNI����Ѐ��RD��Rb _LA`PJͱ��P�pUq|-��#��q�O��XPc�NN�PKET�
��Pq�Uq} h�ARSIZE5p��=���u�S̀OR��F�ORMAT�Pg�C�Oנq�<bEM�d�����UX��,�5p��PLIb�Uq~ � $�pP_SWiI�`��HqAXG�~b�AL_ o�J��A�rB���C�r�D��$EL����C_lі� �� � ���r��J�30 �r��TIA4�Z�5Z�6�rMOM���f��s���pB��ADf��s����PU�NR����s�������P��Rt�� A$PI�&E�kq E�p-~-�-��WC�0$��&��9q�gE��eSPEEDL@G�����Ծ ����)�9����)�8�	)���SAMWPx�p0�1��MOVD� H$_S`Y%nk%_��	1�t�2�t����c��v��8�H�PxIN ����������(�+(+GAMM�<Vu!�$GETHE�U�ٓD5��r
�POLIBRv���I�$HI�_L�ݰpB�&E�(A�.� �&LW�-�&�,�)	6�&�1��f�`j��� ?$PDCK���"ٓ_���r�E� ��b7��a4��a9�� $I��R��`D�c�b~�Ե`L�E�qkq���81��0�q��`Vp�P/a?UR_SCR��A��r��S_SAVEc_D��8Ex�NO5�C��y�6�8@{$E�. {I��G	{I�@�J�KP �q��H� ���x" Mao���s���� d��6W2U�Cqy��9L�0Rt� �k�F� �aE��3�W<�@[�BjQWg@5r�U�R�R���Sc2jQM"��[C�L�W��M)ATr� ?� $PY����g$W`�fNG� O�`�b�b�b #�HЈ��a� ���c��%X�O���Z�e��ހRt� p䠰p�3+zO�O�O�O�O�a:5�_�r� |�E� 8@��>vs�>v��8@_�kwVvy�Eހu%��"rJB�\�P�"tP���PM&�QU5 �� 8*�QCO�U�1��QTH#pH{OL<�QHYS��3ESe�qUE�p.B�Z�O��  q�P����%��UNְ�Q� ��OE��p� �P2�3��AÔ�R�OG�����Q2(�O�}�2������INFO�q� #�e���ڗRȾ�OI��� =(�0SLEQ�с �рi�C�{�D��L���`� OK0r���!E� NU!��A�UTTA�COPY�q� ?��`@ML�NHI�M�X�Cᐛ� Y�_RGADJ�q�i�X�Q��$ഖ�`
��W��P���0���l����EX8�YC0bI�ѪObp�q���n$�_NA9!��������`��� � Q���PORp�A�B�SRV0��)a�Y�DI��T_ ��{��������������5��6��7��8�y���S8BL��m�M�C_F�p��PL9A8An�ȰR��9��р���$iB����d� ,�0FL-`L�C@SYN�[�M��C?��PWRc��L���!�DELA��8Y�5�AD�a��QSwKIP� �Q�Z4�OR`NT�Q ��P_4��ַ@lb Yp������ ����Ƞ��ՠ���������9�1�J2Rܻ L�� 4*�EXs TQ%����(Q�����p�����p���RD�Cf� �`��X9�R�p�����r��~A$RGEAR_� sIOT�2FLG��vi��M%PC��B�U�M_����J2TH�2N'�� 1������G8 T00 I�����MlѺ`I�\8��REFr1�q� l�h��ENA9B{�(cTPE�0� 1���i�m���^QB#���:��"������2�ҙ����������
&�3�Қ7�I�[�m�(��&�4�қ�����������&�5�Ҝ�1�C�U�g�y���&�6�ҝ����������
&�7�Ҟ+=Oa(s�&�8�ҟ������&�SMS�K�q�|��a��E�?AeQREMOT-EF����a@���(Q�IOQ5�I8c(P�POW�0L�� �pZ����#p�%�L��U�"$DS?B_SIGN�1)Q�%���Cl��S23�2��b�iDEVICEUS�,R'R�PARIT��D!O�PBIT`QY�O?WCONTR;�(QX��O'RCU� MDS�UXTASKT3Nx�p[0�$TATU`PK��S�0L�����p_,PC9�$F�REEFROMS8p��%�GET�0��UPD(�A�2U#P|� J��� !)$USA^���6<���ERIO�P@&bpRY�5:"_>@ �qP}1�!�6WRKI�[D���6��aFR�IENDmQ�P$�UFw���0TOO�LFMY�t$L�ENGTH_VT�l�FIR�`-C�RSyEN ;IUFINR:]��RGI�1ӐOAITI��4GXӱlCI�FG2�7G1�0�Ѐ3�B�GPR� A��O_~ +0!�1R�EЀ�E3�e�TCp���Q�AV �G8��"J���u1~! � �J�8�%��%m��5�|0G4�X _0*)�L|�T�3H6��8P���%r4E3GU�W�P�W�R�TD����T���а��Q�Tm�$V 2����1��R�91�8�02�;2/k3�;3�:iva�9=i��aa�^S�jR$V��SBV�EV'�V�B
K�����&c�p���F�"{�@�2q�PS�E��$.rRC���o$AŠFwPR��Gv]U�cS'�� 7�8��E2I�� 0�@qV"`��p�d`���E0��@��=�
B5S!� ��aRg����iR�6�N AX�!�$�A�0L(A���rTHIC�1Y���h��t1TFEI��q�uIOF_CH�3�qI�G�a�pG1bxf����m���S@��_JFf��PR�ֱ�S��~Ԁ�d �$S�z��Z�GROU��̃TOT�t̃DSP�JOG���#��_P��"O������j��&KEP(�IR�����@M�R@�AP��Qn�E^�`�!�[�ScYS6��"[�PGu��BRK�B �.��pIq�p��M���΂�`�AD�!̃9�BSO�C׆�NӕDUM�MY14�p@SV��PDE_OP�#S�FSPD_OVR�=���C���OIR�CNm0�F.�l���OV��SFR��pU���Fn��!#��C8��A�"LCH����FРOV�s0��W�@1M��ĥ:�RO�#ߑr�_�p�� @@��u@VER�ps0OF�Su@CV? �2WD�6���2�ߑj2Y���T�R�!���E_F�DOY�MB_CM4�D�B�BL�b>�f��attV"Q�240/pd��N�Gg�z�AMx�`Z�0���¿_M~���"7����8$CA��7�D����HB�K81��IO�58���QPPA�=��"�M�5�͵���DVC_DBxC~� �3"�Т�!��1��糖�3����pН�*��qU�3��CAB���2VӆPѣIP��c�O���UX�SUBCPU�r	�S�P P� ��90^SQ׹c��."��?$HW_C�Т���S��cA�A�pl$�UNIT��l��A�TTRI"���	�C�YCL��NECA���J�FLTR_2_FI_�G(��9&�1�LP�?�>�_SCmT�CF_��F_�܌6��FS8!����CHA�1�wᇲ�"v�RSD�4"����qv�_T��PRO��,>�� EMy_ܠ��98d��a d��a���DIb0!�RAI�LAC��9RM��L!OÐ C��Q*q��X3q���PR��SQI�pU�Cr�s 	��FUNC��@rRI�N'PѸ0��u��!RA��B ����F��Ğ�WAR~���BLQ����A��������DA����	����LD)0��Q1�q��*q1TI2rQǁv�p$xPRIA1V�"AFB�P�!|�ߠ�<`�R���MO9I��A�DF_&@��l51��LM��FA�@�HRDY�4ORG�6 H���A�0 �MULSE&@"�Q��a� �G�	������$d$�1�$1 ���0���o� xm�EG�̃�`ARހ���09�2o��z�AX]E�ROB�W�A2��_�œSY���t���S�WRI�@rs1��STR��� ��(�E�� 	%1��AB( �/&X�a�ӰOT0^�;	$ߠARY�sf"h���S@	�FI��~*�$LINK����!�a_%#�t%{q�"XYZ828�*�q�#OFF���")�"�(j B�j��4С��n�3FI���%7�q���j���_�J���%��#�QOP�_>$H+5�3�PTB�\1�2C��i�DU��&62�TURN ��2r�5t!}��p��|7FL�`���m�0�%�+*7�	� 1�J. K�M�&82�pQ�2rQ�#�ORQ�� G��-(�+p��z�� �3q�E"��T�GOV�@-A��M*�y�4�E:�E@�FW�J��G ���D��o�*� ��A 7�P��y��E�A�GZU0:ZU�CG�ER���	6�E���B�TA FQ��)4����r'�AXУa2.q�c �W�c�W�c�W�p�Z�0 �Z�0�Z%@�ZK@�Z� �Z
!�V� �Y� 
i�  i� *i� :i� Ji� �Zi� ji� zi�a�iD7EBU{�$v�u���;q��"F7O�n�A!B��6��CV�z� 
fr����uk� �w�!�w�!�w�1�w�1 �w%A�wKA�w��\0���"3LAB"2�|EwЄ�҂�3 &} EERVEN�� � $q�_NmAǁ!_�PO�����` f�M�_MR}A��� d  9T���ERR�����~ TYi��RI�V8"0�S��TOQ�T)P!L��T�ЅL�G�}CJ � p�PqTl X���_V1�bP�Q���#�2�2+������/@��p��5��$W��V���VN�[�$�@�� �S����Q�	EHELL�_CFGN�� 5%�B_BASƴ�SRvp0�K� E�S��Jϐ1a�U%Α2�3�4�U5�6�7�8�RO���� � NL:�3ABn��АACKwv��)�o�pu0iႩ_PU2��COq��OU��P���ӕ�����T=P�_KAR�0&��REm�� P��z QUE٩��@����CSTOPI_ALzs��� �T���� SEM[�w�k��Mw�y�TY��SO`��DI���Є�=��װ_TMK�MA'NRQζ� E���$KEYSWI�TCH��Ѱ��H=E��BEAT��R�EpLE����&�U���Fd�����SO_�HOM� O��REF�@PRi��R� ʞ�C@�O0�p EC�O���� _IOC1M�4M�k�����'�O� D�!ۧH�	U��;�M7��@�3�FORCߣ�� �x��OMq �� @Etxk�U#P�o1B�O�o3B�4�x�NPX_AS� 0ݐADD|��(�$SIZߡ�$VAR�TKIPr�q�G�A(����
�˨r�t�n��SV�XC����FRIF�R��S%�7�xĆ��NFѲEАO�� x�PSIڂTE�C*�%CSGL=�T�"�0&�V�D��>�OSTMT
�o�P\��BW�@?�SHO9Ww��P�SV� K߹� ���A00�0�Q��K���O���P_���i���5��6��U7��8��9��A�� ���6������20��F��
 ����U ���� � ����0�� �J@���:�1G�1T�1a�1�n�1{�1��2��2���2��2��2��2��2�2 �2-�2�:�2G�2T�2a�2�n�2{�2��3��3���3��3��3��3��3�3 �3-�3�:�3G�3T�3a�3�n�3{�3��454���4��4��4��4��4�4 �4-�4�:�4G�4T�4a�4�n�4{�4��555���5��5��5��5��5�5 �5-�5�:�5G�5T�5a�5�n�5{�5��656���6��6��6��6��6�6 �6-�6�:�6G�6T�6a�6�n�6{�6��757���7��7��7��7��7�7 �7-�7�:�7G�7T�7a�7�n�7{�7��K�VP�$�UPD�� � �P���x�YS�LO��� � ���հ�����QTApS�sTƠ��ALU}UL����CU��WFdQ�ID_Lѳ�UHI��ZI�$FILE1_Σ�T�$u�_V;SA��� h��+`?E_BLCK(�8b|g�AhD_CPUQi ��Qi���Sod_R1��ɢR ��
P�W,�d� �aLA��S���c�a�dRUN5��a�d�a�d��5�p�a�d�a�d �T�p�ACC���Xw -$&qLEN~� 3t��&p����Iѱ
�LOW_AXI(�SF1&q�T2mwM��ɢ����I����Q��yTOR.�&p�{DxW��s�LACE����&p�����_MA�uйv�u�w�qTCV�|��wTڱ�;�1�@<ѷt��_��s��J����M����J����u)���u2q2���������s�pJKцV�K~�か��3ՃJ�0���JJ�JJ��AAL������4�5Xr;�N1�B�N��	��tL�p_�k��'*!q���� `5`GROU�PY�ӲB$�NFL�IC�ө�REQUwIREv�EBUV�0"q���кp2���#p�ɖ!qxг�� \^��APPRՐC��ڜp
!�EN�CL9Oz�,�S_M ����A��u
!q��� 䣠MC�r;�Xr|�'_MGц�C��,`p��N��p��BRK��GNOL������Rϰ�_LI��է����JޠѤP��p��p�� �p;��pD��p6�K���8��n�"q���G� ҒMr:ql�<Gqz�PATHv���@����Rx�������pCNR�CA��է�6��IN%rUC�pwQZ�Cd�UM�Yop�����QE:p�Gp������PAYLOA�ͧJ2LHPR_A	NqQ�L�`[�W�K��g���R_F2LS3HRё�LO\�������ACRL�_�����޷C�XrH��P"�$H���FWLEX� qJ%u� :2Dv�p 4�K�GYq�pPbt|F1Kљխ׃�������E��� �/�A�S�e�w����� y���ф���蘏����$J�ÊT���X���� υ ��څ��[���� 
�� �)��;�D�V��h�z�Y�J��� �� �������QIPA�T��ё��EL4� ��ؘJ���ߐJ�E��CTRޱ��T�N��F�ɗHAN/D_VBp�ѹPn`�� $&�F2��K��ШRSW9 qj��� $$M��}�R��E��Uw�H��sA�PH����Q����A���P��A��A�ɫ���j`��D��D�ɫP��G�`1)STЮ�9!��9!N̨DY �`���|�Y�鰋� KыǦ�J�ч�s�U�ХP��&�/�8�A�pJ�S�=��� ;� �t�.R66N�/QAS�YM����Ґ���p�Խ��ٿ_SH�� ���筈4��+�=�O�JV��h�'CI\����_VI�dH|N�u@V_UNI���D���J҅�B�%�B �̦D�ųD�F�̓��� �����*Uc����Y��H�`���XQEN� v�DIɠS�OwT�Y�YP���� ��I�1A �Q�äQ�`Bc�S`� � p�a.a� � ME����R'R�1TkPPT�0) ���Qz�~���0�Xa�	iT@� $�DUMMY1��o$PS_��RF���)$Pf�aLAƏ�YP�jb�S$GLB_T>mU�e��PpQ p���Q� �X	�ɗ`�ST���ߐSBR��M21�_V��8$SV_�ER��OÐ�c�cC)L�`�bA5�O�RTP�T O�P � D� �`OB���LO˰&uq9c�`r�0�SYSqADR��TP�PTCHb �� ,&����W7_NA���tz��9SR���l =��M�u`�y s�u~�s��s�� ���������0�) �T�"�5�~���B�����s�?�?�?DY�XS�CRE)�p�fȐST[�s}�P�!��tX�r _� Aq� T	��`ob���a`�l��Ҥ��g�Zc�O� IS�c���T&Y�UE�T� ��ñjp^`Sq�R�SM_iqmUUNE�XCEPlV֑XPS_�a����޳����޳R�COU�ҒS�o 1�d�UE�t�ҘR�b9�PROG�M� FL�$C�U�`PO?Q�д�I�_�PH�� � �8џ�_HEP������PRY ?���`Ab_�?dGb��O�US�� � @��`v$BUTT��RV`��COLU�M��U3�SERV<x��PANE� qu��P@GEU��<�F���q)$HE�LPB�l2ETER��)_��m�Am��� l���l�0l�0l�0�Q�INf��S@N(0�� ǧ1����ޠo �)�LNkr'� ��`T�_B����$H�b TEX�*��ja>�REL�V��DIP>�P�"�M�M3�?,i�0ð�N�jae���USR�VIEWq� <Ե`�PU�PNFyI� ��FOCUPn��PRIa0m@`�(Q��TRIPzq�m�UNP�T� �f0��mUWARN|lU��SRTOL�u����3�O�3O;RN3�RAU�6�9TK�vw�VI͑�U�� $V�P�ATH��V�CAC�H�LOG�נ�LIM�B���xv���HOST�r!��R��R<�OBOT��s��IM�� gdS )} 2����a���a���VCPU_AVA�ILeb��EX��!W1N��=�>f1?e1L?e1 n�S���P�$BACKLA�S��u�n���p� � fPC�3�@$�TOOL�t$n�_wJMPd� ݽ��U$SS�C6���SHIF ��S�AP`V��tĐG�R+�^P�OSUR�W�P�RADI��P�_ cb���|a�Qzr|��LU�A$OUT?PUT_BMc�J�IM���2��=@zr��wTIL��SCOL���C����ҭ�Һ� ���������o�od�5�?��Ȧ2Ƣ%#*�0�T���vy�DJU2Ѭ�� �WAITU����n����%��NE>u�YB�O� �� c$UPvtfaSB�	wTPE/�NEC�р� �ؐ�`0�R�6�(�Q��� ش�SBL�TM[���q��9p����.p�OP��M�ASf�_DO�r
dATZpD�J����|Zp�DELAYng�JOذ��q�3� ���v0��vx��,d9pY_���	�7"\��Ѽ�rP? N�ZwABC�u� ���c"�ӛ�
X`�$$�C��������!X`N�� � VIRqT���/� ABSf��u�1 �%�� <  QP�/�/
??.?@?R? d?v?�?�?�?�?�?�? �?OO*O<ONO`OrO �O�O�O�O�O�O�O_ _&_8_J_\_n_�_�_ �_�_�_�_�_�_o"o 4oFoXojo|o�o�o�o��o�o�o�o}� ��A�XLMT�s�n�#  �tIN&8qtPREO��+v�upXuLARMRECOV �)xXrzujF �%_�!d ������7�I�[�m�~�,� �/���uNG5� �+	? =#�
ڏ싾� PPLIC5�?��%upՁ�Handling�Tool -� �
V7.70P/�36 ��
]�_3SW2�D�F0j�W� 43Y�J�9�K��7DA7?�����
&�X�e	-�N�one��J������ �T7�	�-rP_�Viu�:6s��UTOz"��,tTy.�HGAPO�N� %��!.�U��Dw 1�y� t��x�����y.�K�Q �1�{  Hp��
����	���uq��"�" �!��Hեw��HTTHKY� �"ٯ����u����� 󿽿Ͽ�����)� ;�M�_�qσϕ��Ϲ� ��������%�7�I� [�m�ߑ��ߵ����� �����!�3�E�W�i� {������������� ��/�A�S�e�w��� ������������ +=Oas��� ����'9 K]o����� ���/#/5/G/Y/ k/}/�/�/�/�/�/�/ �/??1?C?U?g?y? �?�?�?�?�?�?�?	O O-O?OQOcOuO�O�O��O�O�O�O���TO�Ā��DO_CL�EAND���{SNM  ɋ���_�_��_�_o��_DSP�DRYR�_��HI!��]@�_}o�o�o�o �o�o�o�o1CU��MAX �bTQNQS�sqXbTB�o�B�>��PLUGGb�cW\o��PRC4`B�PE]klo^�rO�r�=o��SEGF;�K �+�6��_�_}�����p��ŏ�0�LAPZo m�/��+�=�O�a�s� ��������͟ߟ�6�TOTAL�v�y6�_USENUZ�g�� HXL�NR��RG_�STRING 1�3�
�M�,�S�
��_I�TEM1��  n 󝬯��Я����� *�<�N�`�r�������຿̿޿��I�/O SIGNA�L��Tryout Mode���InpB�Sim�ulated���OutT�OV�ERRW` = 1�00��In c�yclHŕ�Prog Abor^����>�Statu�s��	Heart�beat��MH� Faul����Aler�����'߀9�K�]�o߁ߓߥ� ^S��^Q������ ��,�>�P�b�t�� ������������8(�:���WOR9��� r���L����������� ��*<N`r��������PO�������9 K]o����� ���/#/5/G/Y/pk/}/�/DEV � -�/�/�/??)? ;?M?_?q?�?�?�?�?��?�?�?OO%O7OPALT��^A��8O �O�O�O�O�O�O�O_ _(_:_L_^_p_�_�_p�_�_�_LOGRIxp ��avO�_*o<oNo`o ro�o�o�o�o�o�o�o &8J\n�_*�R�ݦqo��� ���(�:�L�^�p� ��������ʏ܏� �<��PREGbNK� �$�r���������̟ ޟ���&�8�J�\��n�����������$�ARG_r�D ?�	�������  	�$�	[�]����.��SBN�_CONFIG S��L�K�F��CII_SAVE  �k�b���TCELLSET�UP ��%  OME_IO���%MOV_H8��¿ȿREP�|���UTOBACK���V�F�RA:\8� X�8���'`��8�\c�,�INIa@8��^�,�MESS�AGz��������ODE_D��}�C����O� ��,�PAUS�!��� ((O��J�\�F�|�j� �ߎ��߲���������B�0�f�t�%�*TSK  5ݒϕϞ/�UPDT����d�����XSCRD�CFG 1��N� ������� &�8�J�\�n���\�n� ���������"�� F��j|�����/e�2�GROU�N����UP_N5Aܰ��	2���_ED��1
��
� �%-BCKEDT-��}�&�p��Ѳ-2�p�8�/�/�8����g2���E/���/��/~/��ED3n/&/�/J/\.�/"?�/�/ED4?�/?��/\.[?�?5?G?ED5�?n?#O�?\.�?jO�?�?ED6ZOO�O�6O\.�O_}O�OED7�O�Ok_�O\.G_�_!_3_ED8�_�o��]-�_Vo�_�_ECD9Fo�_�o"o]-0�o�oio{oCRoY_ Vh�]1�{� ~LNO_DEL�GE_UNUS�E	LAL_OUT V��WD_ABOR����~�5�ITR_R�TN�ǀH�NON�S)Ю�����CA�M_PARAM �1����
 8�
SONY XC�-56 2345�67890Y ��f�@���?�>W�( А��8��h�х�ڎ��HR�5ǃ��	��R57<0�B�Affފ� �����ڟ�ǟ�"� ��F�X�3�|���i����į!�CE_RIA�_I������Ff��;�Я ����GP 1���s������V�C󠸾����C�O�C ��(��ǀC�8��@��H��CCYX����Ch��p��}x���� C�����Ⱥ��+�=�G���ށ��HE/pON�FIG=�f�G_P_RI 1�B� $r�����������(�~�CHKPAU�S�� 1���� ,wuj�|ߎߠ߲��� ��������0�B�T�@f�x����D�O����T��_MORGRP 2?�� �\�� 	  �,��P�>�t�b���D5�����e�.�?a�a�����K���d��P�V��aÃ-`�/A�

 s�������br&�i��ܦPDB������)
mc:cpmidbg�̼:�~���a����p�U  W �~�c~�d3a� ��d�~���p.{C�eU�/��/��{g�T+/�l/�m{f/�s/i�u/�
DEF 3�(K�)�b buf.txt�/��/��_MC������z/23�����ʇ�Cz  �B�p�B�Z�B��X�B��~C�� Cޢ�D�3�u
q�Dv���D:�"Df���ENNEA�7EV�ߓ=F��pgF=C�Fi��WG���Gp?��G�/�	ބ�	6����4T���(D~��%�/��ʄ3@à1g/  TB�D�V@�2EI�5� F�*� F�G$���F[� GR��kNGl��G����G��&H����G֓�H���߃]��  >�3�3 �ށ� � n^��@߂5Y��Ed��A��=L���<#�
 ��_�*2RSMOFS��.^�9�T1��DE ���l 
 Q�;��P  0_*_>T�EST�"__��R����#o^6C@A�KY��Qo2I��B�0�� �C�q�eT�pFPROG� %�S�o�gI��qRu����dKEY?_TBL  6���y� �	
��� !"#$%�&'()*+,-�./01��:;<=>?@ABC� �GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~����������������������������������������������������������������������������q�������������������������������������������������������������Eъ`L�CK�l���`�`ST�AT�c_AUT/O_DO��O��INDT_ENB�;���R�QY�K�T2����STO�~���TRL�`LETE��ފ_SCRE�EN j�kcsc 	�U�πMMENU 1�i  < �l�ol�K�u���FS ����柽�ϟ��� R�)�;�a���q���Я �����ݯ��N�%� 7���[�m�������ɿ �ٿ�8��!�n�E� W�}϶ύϟ������� "����1�j�A�Sߠ� w߉��߭߿������ �T�+�=��a�s�� ���������>�� '�M���]�o������� ������:#p�)+�_MANUAyLӏ��DBCOu��RIG�$�DBN_UMLIM�,1�e
�PXWOR/K 1k�_�-<_N`r�TB_�  m��Y0|�_AWAY�%�1G�@b=�P��_AL� =���Y�Ҁ��`�_�  1}!�[ , 

�:&d2/o/�&�M�t�IZP�@P�#OoNTIM��d���&�
�e#M?OTNEND�o$�RECORD 1�'kU2)?�!�O�?1-?&k�k?}?�? �?88�?�???�?c?O *O<O�?�?rO�?�OO �O�O�O�O�O_�O8_ �O\_n_�_�__�_%_ �_I_�_o"o4o�_Xo �_|o�_�o�o�o�oEo �oio�oBTfx �o��/��� ��>�)�7�t�� p u�����-��͏ۏ� ����N�`�Ϗ��o�� ��)�;������8� ��\�˟ݟ����;�Q� گI���m��4�F�X���TOLERE�NC�B�	"�L��Ͱ CS_CF�G ( +x'd�MC:\��L%04d.CSVY�� cֿx#A ��CH�z _/x.��G��},��RC_O_UT )�- �z/��SGN *���"��#��17-JUL-25 20:52���27-MA}Y��14:38��]� Z�t������x.����pa��m��PJP���k�VERSIO�N ��V�2.0.11~+E�FLOGIC 1�+� 	d���ٓ��p�PROG_ENB�2��WULS�' �p�_WRSTJN� ���"�EMO_O�PT_SL ?	��]�
 	Rg575x#?�74D�56E�7E�50i�dԂo�2E�d��j�"�TO  .����k�[V_� EX�d�%� �PATH A��A\��M�_��~+ICT�F��, '�`��eg��}�STBF_TTS�(�	��E��`���� MAU���ߧ"MSW��-D )��},t���.�!��]l�R�v������4SBL__FAULy�/�|�#GPMSK��^�"TDIA��0����`���!1�234567890xS�l�P��� ��//%/7/I/[/ m//�/�/�/�/�/LZ0PV �� �/�2?X?j?|? �?�?�?�?�?�?�?O�O0OBOTOfO8<x�U3MP$�I� �A�TR>�O�@PM�E���OY_TEM=P��È�3��4󜐰�DUNI	�w�Y�N_BRK 1���x�EMGDI_�STA	��GUNC�2_SCR 27[��_�_�_�_�& �_�_o o2or�nSUQ13y_+?|o�o�o�o�lRTd47[� Q��o�o���_>Pb t������� ��(�:�L�^�p��� ���� ?Ǐُ�0�,p ��+�=�O�a�s��� ������͟ߟ��� '�9�K�]�o������� ��ɯ�����#�5� G�Y�k�}�������ſ ׿�����1�C�U� g�yϋϝ�ׯ������ ��	��-�?�Q�c�u� �ߙ߽߫�������� �)�;�M�_�q��� �����������%� 7�I�[�m�������� ��������!3E W��{����� ��/ASe w������� //+/=/wa/s/�/ �/�/�/�/�/�/?? '?9?K?]?o?�?�?�? �?�?�?�?�?OK/5O GOYOkO}O�O�O�O�O �O�O�O__1_C_U_�g_y_�_�_�_�gETMODE 15'E�fa t�|�_GgRROR_PROG %�Z�%���HogTAB_LE  �[1O��o�o�o�ZRRSE�V_NUM �R?  ��Q�`�a_AUTO_ENB  u�SZdw_NO�a 6�[��Q�b  *�*6p�6p�6p�6p�`�+5pOastHI�S�cXa�P{_AL�M 17�[ �2��6|6`+t�@��&�8�J�x_�b.p  �[4q�R����PTCP_VE/R !�Z!6oZ��$EXTLOG_7REQ�v�y��SIZ�܄TOL�  XaDz�r��=#�
ނ_B�WDo�%��fQ���_�DI?� 8'E�t�TXa b[�ST�EPg�y��P��OP�_DO�v$v`F�EATURE �9'EQ��Q�Handling�Tool � D�ER Eng�lish Dictionary��7 (RAA� Vis"� Ma�ster���
�TE0�nalog� I/O��p1�
0�uto S�oftware �Updateb� �"/�k�matic Backup
��d
!��g�round Ed�itB�  25L�Camer�aT�FX� "Loμ�ellT��L,� P��omm9�syhۡ�h600��scou���uct���p�pane� D�IF���tyle selectѡ;- /�Con��9�?onitor���Hd�tr�Rel�iabT�ϣ(R-�Diagno�s��Q�	�H�Dua�l Check �Safety U�IFc�Enhan�ced Rob �Serv��q ��v	ԸUser� Fr���T_i��xt. DIO� f�fi�� )�\��endܰErrzu�L��  prנ�*�rO�� @���E�NFCTN /Menuİv�����.fd`�TP I�n?�faco�  �
E�G��p;�k Excذg�C���High-Spe�ܰSki��  P�ar+�H���mm�unic��onsn��\ap��urf��?�X�t\h8�U���connZ�2�Т !�Incr���str)�8��M�-6�KAREL Cmd. L���ua��}��B�Ru�n-Ti�EnvB�(<�@�I�<�+��]s��S/W�"H��Licens�e���� ad���o�gBook(Sy�>�m)	���"MACROs,�¿/Offse\�fĜ���H�!�Y�M1��MechSto?p ProtZ�3�o 5
�Mi4��Shif\��B6S�MixܰQ�����H�Mode S�witchY�MoTk���.�� ��Mt�Q�g�� �5��ulti-T�������)�Posj�Regyi>���  ! �}PA�t Fun1מ�6iB/��R�NCum�Y�3�G�P/�|�� Adju���	�/2HS�)� yo(�8�tatu����AD ��RDM�ޱot�scove&� #e�v�㱗���uest 86�7.��o�\���SNPX b��Y��Þ)�Libr%�
�r't I���� "���Ҫ�.S�o� ��s in VCCM����� j������㣀/I�� 71�0�TMILIB�X����g�Accܨ���C/2�TP�TX�� �Teln���Y@����K�PC�Unexce{ptܰmotn��� ������\m725����w�5����  h640S?P CSXC�i �� j*�� RIN��We���50,���vrl�زme�n" ��fiP-�a����P��Grid�{�play F �O/��? ��ELR�;�|�20��OR�DK�sciiw�l�oad�41d�s�t�Patd��C�ycT�h���ori�ɰ:�7c Data&� qu6�2�0�*�p������FRL�amc�K�HMI �De��(����k�P�C�φ�Passwword�644���Sp�����D#YELLOW BO�	�?1�Arc%�vi�su����#ti�OpX�^�! 2��aO��po�� t��ֶT11o�����HT���xy�	�   $�t۠ig��10�Ơ 41\+�JP�N ARCPSU� PR+�8b!O�L0Sup�2fi�l� �!��E@-�;�croc�82��v���n$ 12jSS0]e4�tex-� I��7�So��tf�ss�ag�� e��У�P���,��� "Tc VGirt��v�!�����dpn�
�J3ނSHADf0MO�VE T�MOS� O TԠg�et_var fails l�>PU�~1E���� Hol�d Bus %�h���VIS UPD�ATE IRTO?RCHMA A�{��vYWELDTV S� ]�DtS: R7[41��ouiPb}��y��BACKGR�OUND EDI�T "RC$REPT�CD CAN C�RASH FRV�R 62z1�SCr}a��s 2-D���r ) "��$F�NO NOT R�E��RED �` �m ��JO� Q�UICKaPOP �FLEN m41�S�Loc��gRTI�MQ%�#�FPLNs: FG��pl m��r`�MD DEV�ICE ASSE�RT WIT P�CV;PB�AN#aA�CCESS M �.pc��Jo��Q�ui±�Kbldm�gUSB$ ��t & remov��� Pg�SMB N�UL� ;a|�FIX���C��ACHIN�,QOL�`MO O�PT ՠa��PP�OST0�WDU �C�wQAdd�`aYd���0io�2��k$P�`W\0.$0`�O�IN&�P:f�ix CPMO-�046 issu5eC�J/aO-�0�r7130Т- ��vR�SET VARIABLES-P{��R�3D m��vie�w d��M��&�e�a���b��of �FD�5P:N@x �OS-1y0`�h isc���t��s t�3lo��7 WA�PZ��3 CNT0 T��/"�ImR�)�c�a �Pu��POT�:Whenapew�B�STY E�{1t���ptKQdo G�ET_�p �p��V�MGR LOl�REAd0C~QW�~1��(�l�s�gD�ECT�pLpING IMPR�DR(p+PB�PROGRAM�E�RIPE:STA�RTU� AIN-�;�ӠM/ASCIyIzPÂOF Lq��DPTTB: Nv�pML$me P����`:x�mo&�a�llW`!�ӤTorBc�A�U�HC�iLp�Ըth�`n�@ c�h��/GEA�!�toyu͐�RCal���k�Sign`� N�D�ԗThresh�123��`��09p : MSG_P��+0er  �Q�Aܠzeron��0� H85��RImlA�n�2D��rc�0�I��OMEa`�pO�NaP5�  נSRGEG:FF-Д� ]�|'���KANJI���n��J��c�0asn� d�!OA imm�c �INISITALIZATI�����~1wem����d}r+� LB A�U�Wqminim�r�ec[�c!�R���m>$�ro -1>ѮS�ܰir��@ұJ�1pdETw�� 5`?�I��ow u��< se� 1lc��YbPM ���p�Q���R`vR&��lu\�3�Re 0��4q�q1#���m <a�arn��ঁ?Box fo��*PORWRI�PW�S���v�09 F�pup~�de-rel2 �d�p� j��`━b�etwe��IND� Q���igE s�nap|�us��s�po TME��T�PD#�DO�p#aH�ANDL 1\kP�`vR��ȀD�ny��S�v�Yopera�bil� �T*�: IH � l\p��Vq�Hb�R�< p�a*�c&2�O�`FA,�.�-QV�7. f.v��G-T�pi�s��� �ɠtmLine-Remark ^�� RM-�` W��#SPATH SA�+PLOOS UIqFc�+5f fig�pGGLA����Vrp�������U�0ther|�V� Trac��"�tW�\b�s7��d��t�� n�@  ����3:���dK�y���it k8�d�P;ayR![2]�ü�1: g��s��d�ow�XQ��0IS��q�qEMCHK ?EXCE C���OMF +�Xah�� 35\k��)���QBt���'b���2[�c���e �`k�<�S�� BUGr�:�cD$`PETp����f�c4��0XPAwNSI��DIG���@OoPmetTCC�RG EN��CEOMENT�A M̀�K {�`H GU�NCHG �`� ECXT�P�2�bQS��93 wP8�x�OR�YLEAKq  �H5gyq�PLC �WRDN R �O9 /u�QSPE=p��G*�V ��$�t�n720\3pGRI��A�rT�PMC� ETH��pSU<7p�`  j5/n�/PENS�PN,���*P ont�`BR�OW�`!sRMV 7ADDz CN q�DC���PT3 A�LA2@ ���pSV�GN EARLY8�R��ŰH57�Ga�JLAYҀE 5(@M�PPD�p*@�H�S I`P�OGUCH8���V�F�q��comH�x ��E�RROR� DE �nJ��RO�CUSRS8pI��N4<q�-158n7�ORSR xP#aUp�P��Rqy�T�Fz��;�pk��t�� g�Ղ�B�SY RwUNN�  a�`��BRKCT�!RyO�p3@ \apS�Ƣ�AXxP���h8x+ q��ISSUrp} sPX�PTSI��K1M10_�IP�SAFETY Ck�ECK[��Á�������<#X�� �T�WD2�@�@�IN=V��D ZOp�5�X��t�DUALy� "M6�0�"r�F#�E��dPdNDEX F�t*UF�"Pʀ�0s�FRVO117 �A�PT6�KtqFA}LPTP2477D�6_�P�!;HIG�� CC�t;SNPX� MM��tq�d~�Vq�q#�
"��DETEC�Tq*@RRU�qA�P�5p
�9 y�)<9���7�T��Pds� �k�	���!Q����� t\4A�;A0�27 "Ke@" 8@HI��qXF8@4@H�PRDC"�
�aMB8@�IXF�b���zOX@8@����a�G}E�B�Ccsc�r�J8@�Ndctrld.�A�NZE�A5�I�Q��!�`�Df8@\�`m�878�Q-;� ��� rm`�
���PR̠78�@RaI8@0q�Q (~\�Mp��0t��!{B8@\PtQ<OX�St0�3hB�3nO�Vtp�A�@L�CF�L��� �Rplcf���J8@�WTa�mai�E8@mubov2_miTA�O�S8@U`�T[tT�AqPr674�xSShape G�en��8@j�I�[R��`�@8@T����%q 1(u8@��II�^�Q�~C�a�[8@;Ynrsg:0�4� � 4�CtMSr68@�r5hB5�z�Vnretsp "�r�Po�wng0bGCRE�Ka�ޠ��DAT�E�k�cr�eat.�q�M�a��oksqgtpadx1P��(�tputZj@�{�������܆28@`����Q����sl�ov��� �hexH��TB�8�ď�keyH�8@�pmZb�NR�1u7A+�nrgc8@UQ��pp�bUZ�dp0aj�921xSpl.Collأcq�\A��R1Nq�UA� (J�8@ip�_�WA��_�Y���a7hB7�ͦtp~[� "TCLS9o<Kb��clskyh[:��s�pkckZd� ��$�TQ���dA�rx��710a- KAR�EL Use S=p�FCTN9�a�a7l�0s0a�� (�� �a��~C8@��MI��c�8hB8"   ��8@ v	��v	   lomatea99�q�M����E�mcclm5�CLM;�� �j̕�E�et���aLM�	�h�yasp,���mc_mot�B�N��`8@H����Q��su'���Q�ȕ�䅮���jo�i#�ߕ��A_loqg�Z���trc�B����ve�ϓ�v��Q�WX��6�finde�rxSCenter� F1�lSw520���ha6rX� (<�r1,�Q�Ձfi�Q � NH0�I�ۡ���A8@uL���tq�a "FN�DRVϳ���etgwuid�UID�C 8@���������TA@�nuf;��P���ƞC�B��_z�Ӡo��q�G������l���fn�drTY��2䁴tcyp"�,qCP MF�:}38@517��6s38�E��gf6�� (��K��Q��-�X��A&�tm6�P�İ ��Q���	�͘���tm�Ĵ�b8@e0j��TAiex��aP��Aa�ذ�cprm�A��l�_vars��
��dwc7 TS0��/�6��ma7AF��Group| sk� Exchang�J 8@�VMASK �H5�0H593 MH0aH5@� 6� +58�!9�!8\�!%4�!2���"(�/�@�;OMI� `@a0hB�0�ՁU4U1#SK (x2�Q�0I�h��)��mq�bWzR�DisplayImQ@QvJ40�Q8aJ�!(P��;� 0a��0�Ϙ� 40;�qvl "DQVL�D쌞�qvBXa`�uGHq��OsC��avrdq8�O�xEsim�K40FsJst]��uDdX@TRgOyB�Bv40)�wA�~���E�Easy �Normal U?til(in�K�11 J553m��0b2v�Q(lV40xU)���������k98�6#8Uϕ�|�rP "NOR��dw d.a}oKksu�O�W���O�Y�W`�j0�6�H� mOenuuyP6�M�`�wRX�R577V�9{0 �RJ989}��49b\�`(�fity�����e�<?L��Vsmh`��8�� C0�Sv�q�8����w�pn "MHMN<��ޣx�Ay`�o�3@�u�`f�І�x�t���tRzQ��LV��vP�tm���|I�1{oPx ��2|���I�3I/B�ogdstǏًmn吼���}ensu_�L<���h!!��Rt��?huserp��0���ʐcM�_l�xP�oxe��рpoper��|��xdetbo/� l>�x���Ps$p�`����OPydspweAb͓��z'R��u�Rr101&S՟{t�`12�Z4�30���D���`4�
�4�5���KQ�m[T��dUCal G40`�Q)p40}������9;��DA��� v	LATAu�mpd�\bbk9�68��68c�fb\l�41969y�9�|��D���bd� "B�BOXêM��sc�hed����m�se�tuM:�����ff ���40��n�41�ϒ�40q�col��|�1�cxc�ؘ���li�� X�0���j��&�8�4 �<�ro5�TP E��#��ryK42�r��;�(T+Q �Rec'�ʈ1Iw�84������Ak971���71�;���parecjo��QNS��[T���dXrai=l| nagek�M �,QT2 *� (�ĜR%<x�80!�bh��p��4��4��yDgl�paxrm?r "XRM�g�l�brf{���n����kl��9turbs�p��㧑- �l0195	�g�625C�M h�+���)89��	+��B6��o�ҹ���x�7�q40����pd "TSPD�=<��tsgl��l��:dQ���8Bct���K�vrE�aܮ�����  c�!���21�`�( AAVM l�2�0 �@fd �TUP him �(J545 �l)�`8 616 �%�VCAM ���CLIO �(�0:�5&  {(F\ MSC �R�t"PBsSTY9L�D!28 :2\ �NRE F2h SC�H6pDCS�U tpsh ?ORSR �rD!�04�SEIO�C& \fxh 54�2 LEX"� E�SETn�8!H ��s�h8 7H �M'ASK�Ø"7>���OCO*`x�!03P"6�!/400:66$ �G639.6[8LCH�!6OPLGR703�
5MHCR��0CЄ (! �06�A.f�8!54
��00DSWb 588�180 ��h!37 88 (%D�"02C24���2'7 q9�25��2�-6�05��9P�RST bBFRDMES�!zB��930 _ NB�A  6� HLBo 3 (~!SM�@� Con� SPV3C �8!20z���TCP aram�\TMIL �A��@PACETP�TX �@p TE�LN 96��29^�%UECK��r UFRM et��P!OR ORP IP�L%CSXC�0j��1CVVF l �FQHTTP satA")�I#� CGHP�8ZIGUI��0�hPPGS T�ool� H8�@d�jZ��!@�h!63��%�@32Q\�31 �B�h!96�%R65�1�Rs�!53 T7FAD�R41�8"[1 ��oo�"9��41775�"/@�P�VCTO�@�U�!s�h!80�%PRXY<�R�!770 �b8 ?885 ol3P� L� аdi� �`ڳ�h LCP{Q� TSS �b�26:����@�CPE �HT@V�RC~�tQNL <��@002 %��b�	0dis� �`7 `<��a\0�T�`1 �`{en�b4 652�`)FU02Q0Πo`dp�Ptu�r4 $�r5N��RU0p@n�se�QJp1 AP�FI[ Jp3�g34>�g40 alxrlE1t44w46� ts U0  7v�0�O��r5�e�p7 po "sw�a61:���r4��r5 QpwGr`�$�p8R�"sP`�tQ�b�36w77��w8`�v83���r8��&:��pOq8�8 "/rkey8�9F��a;90�91 p�#@���� �D095�g9-7*pur�A1@d����P|P�q1�0Qpl�Sq1p#4��]a!s1&@sl༂8�Ӽ�$\1�d1�`��v�@�{�14p�ae��5 �h2��`�6ޣ��7�f1p@��d�YpCqd�ـd�1�`uq��� BCu1< Oq� ��7ReU1$ �u1�Pϱ� ܺ�@- WQ158 ase C���9 B��60 8�2ń�p���4 (Wai��`吢!��i7E��8�EU1P`�ro9�<�1��<�2 ��<�	0��T��l��5J�l��cC���9�%�MCR��P�2��`�Q2@967��Q��8��9Z�2�TPB���P�2P7UA5@�o���
�5�`U���3 w���?AH�E�1��c�qAwl���A�1��512 f��1�u5Р���a5p$��56�+a��bQ5h��Ұ�1 @���pp�b[�538� xaB��|p�4�2��11/q5�p�4U5�P16 (߲�Pz��0��8�P����$�p�e5`�e5(�/�P`bbf>�X��$Z��U�5d�\� ~X�7 	  �ÿ8 k_kv��7s9 s�82 &�H5��E6���p����Ah���ñ���3J"ܫ`��4 3Ȥ59Jѧ6�0t���8��q6D0$�$�4 7���!���<�j670\tchk<�Ps0��<�B<�90��7�H<���<�\K�<�q�� ��A�C<���q�<����<�t��sg<�lc$���FA<�H��<�`��<Я���<�hk�� <Щ�B<е�o�<����<��K�<�dflr0��<Ш��� ��oҠ`���D�;�<�gEvam����B<г�o������<а�KЀ�creexl����P��<���|���j6<�s��prs.`���\���<�7������f�sgn��P�b�t�at��<�L��1B >!�svsch/  �Servo S���ule>�SVS��44�1u�_<���� (����ched���,��~��A\�� �� B���B�qA�����cj�� � 5��1<���Ә�p�css "ACS<� &(��6� �����c el���Q���~��torchms�n<�- T�Ma`�x����09 J5;�598 J681
s�7� 8��b���<Чa����te,�s�����/�E��s m��ARC.�� 1q�4�!=��C�tc�pA�@t�L��f� F����7#�2x�SE�r����UtmS�0960'���RC���`���� p��96G0= '��"H5W�� ��L���\f��� �PATb���`!40U�#!Stmt��E ��� �pMA��!p��z�2?�inA_<�X��r�X e/	cW����V���чetdl�vߏ\oveto���܏��mmonitr�0\��|#�0st��?.6a��PP����! Q�!y`�`am9e �Arol�c�43�0 �p��6��01� 25��  �<� ?v	�v	�A@�818\n; <s��I�B�2�pMPTP�"��C�1mocol��,��CT�v�'!� 0�A���8P53��y`_Touchs�s�`��<��J5���� �`mP����n[PQ �a,�E�a��IP&
&�Pth�A<�KF#R��m;�Qetth�TGHSR'�q-�Rt��o "PGIO�#�!$s�ISwka�"W�K��!�MHqH+54��5w5n/�Sm/��@ 7�*�da���8`!w/Ac��tsnf Tk�/�#gb��a��u`��^m�`u ��Zӭ�ܱQp�є� #���Ka<��M��t5QtZ�a<��dFS�5GK����G�1or��dW��64��tPx� ��P ����x,�� ?$���P<�Z4e7�g "SVGN.o�x�copy "C�O;�Wj$�O�A�9� "FSG�ѧ�%7���_��f� wQSW�F*!"(�sgatu`ɀ���_
��tp_�TPDo��9�7�9�#dߎ?���h�G�AT���!#��  �Гf�` ��" /� �w�Z� �b?6?�  ����� ���E ���M� �chrT� �K6K� �sms� �o6��~��gtdmen?3� �?��� ���mkpdtd2 ���, ���pdQ�X� ����� ����mvbkup.� �[�C�С��mku�no��prp���m�kl �4��s �n�iU��� �ldvrw���glg�4�� �p�棑��aut7�.pб�旐 �ַ������su3� �Ǜ�  �Ƿ� ���\ �6�b2X� ��&�� ���<��A4�  ��B�   946"� ��fB� �t\pa�ic\p4k94�7 ���F#���� �i�ctas���pa`���cc:�<��o������gen�� � $��F�lnp � �����stf@��1��wb�O�c��Ջ�`��߄�vri�ߢ�а�-T�� ���p�flowl� OPAc��ow���R50qtS �#T� (A��4�#���pѣV�cu3�QF�� ��SI�ac����4�6����s&��pa���!!���� ���55 �b �o)�p���0娿>
�afcal3�P߁ ��f��}���`�f��m	߳�p�d�m�/���a/��$C`ѷ��� �! track�\P� 0�ine/R?ail Tr�]T�J�69W�T  (L ��8(`љT.�`�%���D��P0� (��8�48��_ɛ�⇒A4����� �3�b13���alV@ ��NTf���%��Ii�n]0m���aen ������&?5�c@Itst3@��$� ���`�,R9�%����0氱%��pop_eners-OW �dDev��F�M�6 W���|A�Pc"�l!esv� �,��R��V$��Q���U<�V$ �k9j �6��# ������%paop/!OP�NU�V ��2celL��8g_��/�6��tscG��$���V!�3� 5vro!p�ߡ�7`�n(`� V"2D�a V'O$:S|9��� PumpE� �jQ�@�" ��!
��@бMSC#�@��)P��A�C�`��� � �v���� \mhplug�@g�"7Pb��uK")㠱io7��CJ0��E�LIOj q1g 7A93շ��5 q9 t����4.rb ST��R��CP�J989�P�LSQE�' �e C3Q(P �/Ov���o�P�� ? I1�R���5�5��f�I1`�tcm;io��MIO������Utco1"CL0�1V �cBK`io"��uM?���Sl�I0�ߢ�Eg �o���f �1tI4\onfdtI����e%�p27�Int�e�TB CoMo�o1E�R�(do5�54 (;r>Ex,p��nR##ipc�/L>��qp5���
oQ é�1�p����7/o��j�ra�pd�CDV�_��rP�֮��qp2c�nd��s �p��a �o�r`҄�S��"�c�1a�c���2kIԿ?A�pcrt���or0�qd#��"���3p+�཈D��Џ��vr2k�0���AG�.+�η�cho�;�uCp��(� �uV630� fwe P�mී�@���,`��TX�� ��d�chp "_��(	�3�����8����\p3�v����ш�9�3�1 ������low�[ͧ���chk���㳦s��s?Ө0�i�1h���2��i�w����s?1*�-0	�:�O��vr����৓0�'���PFRA�PWat?1rne@E�P�sp�& ac5� \_A�rbo#�,�a ��g��������Q=s<�ICSP+ �9_����� �q�F�A9PH51IQK93 7��HX6hQ�]PVR`S5��fPR6� iQWPR� (P^!am S�u�"��A�I0�tpprg��0���`h�@2atk932�!��E�^�^�asc "8�C��S>i�atp�"�d��@1I�
g�dsb�lfltJA�Qsable Fau�P{C!��EV0ex/!?DSB (DC��t�$�p��X 7�  �� 5��Q�t3*�~l���td9� "!0%�(5��sb9኏���\	�6#���@5��p$D@550-Ad�just PointO"tVJ�Rs�z�@䐄��!�X_�Yj�^�0\sg��4�߼}7y�\ada�"�ADJ���j�Qe�tsha<�SHAqP�sŭ'jpo�r 4�t�!��$ ��C�|�	Tk!bRPK�AR/Qiagno�stì!O!vV6�6 J`ew0�(��L���/�&krlde� ��PP���h�U b���r3�Pp<?q��DBG2C��� �X�o�1U��� ��WT`�@ip�JCM�aipper� Opv`1Se}78 (MH GF�  ;":�&##�� a�xX�֕$��388C�P����#��9.�9C�H�g##PPk�Q��8�! �_"$�"��=0%�P��A  $��_�#%0AQ�C~2� Mat.Han�dlE��!= &�pq MPLGET�0�1(�3�Tt&P�Sٰ'�B �1��B0����&p��H ��PP �'p��@�C7�PP	�TG�tD5�}m��q�Afhnd "�F_R  ���|��PP	   xT�?Q���P(Pa��TAo�����?�pmp�aO��JP ak92�5��2`@O�JRp�sQ`B2�unLHP�Tgse�GSo1�O�W�QT��v !�R�P�tp~���JRdmoan.�@��V�!ns�hYvr�QJ�g�Q�o��jY�HS~7sl�f .��pen�PDnR(R8&���ɐ823'�� ٔq���g� ���� 1��� S�� ? �c\sltQ�!|QE�P��a�r�tPg��P�� �v��"SEDG8�s0�qtdgY T��� �vP`ho�s`<`����qc�`g
�e` op�w�a@o"�ile6�H�e�ȅnR�� x�e! j517�>Ճ��J%��e�`��Q4��Q&�L�!F�J�=�o�5�z/l17���_�œ���`C0C�  ���LANG j��A���8�����gad��X�#�jp�.�0�4�Ē�ib���s�Ƒpa����&���j539.f��,Ru� Env
������3H�z�J9�����@h�Ф
Ҕ���2�a2���� (KL�n-TimФ�⠤���p�3�TS����\�kl�UTIL"�o���x�r "QM�Gl��!������1� "��S�T3�\kcmno��SФT2����ut�.�lrgeadc�}�exY�(ܤ�r��\��l��Ф�w�3��2C�*� - �C�D�E!Ĥ� .��C� R CV̴�Ҁ�C\p�Р���pďtbox��.�@�c�ycsL�:�RBT�E�veriOPTNE���;ӕ�k��e�ߦ�a�ߦ�hg��ߥ�DPN��gp�.v��r�ptl�it��0�4��te\cy����tmnu3`�r�����5UPDT��������駣��i�te �� swt�o�,���oolB �F"�Y���Q��(q��gr3��䪒��"�䴁w������߳��s��������������lS���bx " O�� ����l����0P���A�l\t�� ���������	�Colr�e!��R C��r��&r �m;`��Chang�Lq�T1 �rcm3�"��
�� 6���"����sP70���"��22!2��2D4�57�� CCF�M�H��accd	a��Q�c' ��K�@�0���K!����mo! ���,$Á��!"
 ����/�/����	Y�`,$��)�,$sk����m rC%tS1,$+�x��k1�%unc.,$poñ�1��sub��p����1��cce�5 /!&��-/?-W/i&vs�}/�%#�#�/�.@C��/� C%
�@? U ��&+��F:qt�
pD�Ѓ D	 � U�:7�Dxmov.�P��DPvc5Q.�tfr@PeC_UY?geobdtg_y[�tu���P���PTUt$�P�Sx�_�^z�_�\gvar�_�\xy�_.�[pcl`c�P���P�Ue�Pgripssuaoskuti��|�ovfinfpo}��o�j�b�P���Qud�\�aX��Pc�\Rrp��Qnƅ�P�v�P)tm�#qƆ�P�v�a+rog��a��\Q�?a+rpal?a{�{spa���P �u�Q�t�_TZp�0�osipkag3r�ovlclay(�:�t�pT�d�pu?a�c�A������KtKa�P��r��qTf|rdm���{rin#r���s � �2���|s�Pd�&v�tv��v�h�0���ystn* џ�yt'�1�p��D�p�uϑ�#�ul�@o�W6�2�siupdl�]�o�#vr�on��`1L�zp�`\�r���il3F$|l4��ǉ#q54�FyB�Տg{�`���{w�cmס���wxfe�r�UYtlk2pyp߿UYconv���sicnv�Qʯxaqg��H�Z�lct`a�o�=�p��׭nit�0믁�3������ � �� v�	�v	$��a�lϑpm�r&�B�e Wa���f�%���� ��I��߬�u�ͬ�Ka�mT�f���c��w��roǁ#�5�����?� sm��y�a��y넑 ������`����͐ϑ��p��m�Wa�1� ��A�6�S�e�X��� ��\Q}����������� ĥw߉�西߭���� ��#q0��rs�ew�@��1�a��z긱n@��.�۲;�d�������  � A�d	T$�1 pc! P��e �e� 	lf@C�@��s/�  ?�����8�� �������re�g.�C=��o�99 ~@�����$FEAT_INDEX  z ��e�� ILECOM�P :���1!!z$#�SETUP2 �;1%;"� � N f!$#_AP2BCK 1<1)?  �)��/��/  %�/�/e 4 �/�/>%�/$?�/H? �/U?~??�?1?�?�? g?�?�? O2O�?VO�? zO�OO�O?O�OcO�O 
_�O._�OR_d_�O�_ _�_�_M_�_q_oo �_<o�_`o�_mo�o%o �oIo�o�oo�o8 J�on�o��3� W�{�"��F�� j�|����/�ď֏e� �����0���T��x� �����=�ҟa���� ��,���P�b�񟆯� ����K��o����� :�ɯ^�����#��� G�ܿ�}�ϡ�6�H� ׿l�����ϝ���@)�t Px/ 2� �*.VR��߅�*�@߂�F�j�T���PCrߛ߅�FR6:����V���z�T �!���K� x��q�S�*.F�D���	�Ӑ���^�<���STM ���'���S���i�Pendant �PanelS���H I���9���U�������GIF0;���8�����JPG���;��]oR�
A�RGNAME.D)Ty�>�\"���Rc	PA�NEL1Y�%@>��e�w��2��A/�//���/�3 _/�/��/p/�/?�4�/I?�7?�/?�?�TPEINS.gXML�?>:\�?�t?�1Custom� Toolbar��?Q�PASSW�ORDg?w�FR�S:\:O�? %�Password Config{O R��OSO�O�O��_�O B_T_�Ox__�_�_=_ �_a_�_�_�_,o�_Po �_Io�oo�o9o�o�o oo�o(:�o^�o �#�G�k� ��6��Z�l���� ���ƏU��y���� ��D�ӏh���a���-� Q���������@� R��v����)�;�Я _������*���N�ݯ r������7�̿޿m� ϑ�&ϵ�ǿ\�뿀� �y϶�E���i���� ��4���X�j��ώ�� ��A�S���w���� B���f��ߊ��+��� O���������>��� ��t����'�����]� ����(��L��p ��5�Yk  �$�Z�~ ��C�g�/� 2/�V/���//�/ ?/�/�/u/
?�/.?@? �/d?�/�?�?)?�?M? �?q?�?O�?<O�?5O rOO�O%O�O�O[O�O O_&_�OJ_�On_�O _�_3_�_W_�_�_�_ "o�_FoXo�_|oo�o��o�`�$FILE�_DGBCK 1�<���`��� ( ��)
SUMMAR�Y.DG�oblM�D:�o*n`D�iag Summ�ary+8j
CONSLOG q�n�=qConsole log��7kpMEMCH�ECK��2���qMemory �Data3�;g� �{)�HADO�W(�����C�S�hadow Ch�anges���c-���)	FTP������=��qm�ment TBD�;�;g0<�)ETHERNET0��`n�q~���=qEthernet �p�figurati�on��B`%�DCSVRF/��'�@�C��%� verify allC�ޑc1p� �DI�FF8��0�ůD�{%Z�diffǯ{��q�1������J�� X�q�|�	�CHGD�&�8��ͿD�ܯ�����2pĿ����R� `�yτ�GD�.�@����D�����FY3p�ϳ���Z� h��ߌ�GD$�6�H����D�����UP?DATES.$�
�~ckFRS:\"��c�>qUpdates Listc��`{PSRBWLD'.CM��blN���e��pPS_ROBOWEL\�6o+�=� loa��o����&���J� ��n�����9��J o���"��X� |#�G�k� d�0�T��� /�C/U/�y//�/ �/>/�/b/�/�/�/-? �/Q?�/b?�??�?:? �?�?p?O�?)O;O�? _O�?�OO|O�OHO�O lO�O_�O7_�O[_m_ �O�_ _�_�_V_�_z_ o�_oEo�_io�_zo �o.o�oRo�o�o�o �oAS�ow�* ��`���+�� O��s������8�͏ ߏn����'��� �]� 쏁������F�۟j� �����5�ğY�k��� �����B����x������C�үg�v��$�FILE_N�PR�]���Y�������MDONLY 1<��~U� 
 �� ۿ(���L��5���Y� �}Ϗ�ϳ�B����� x�ߜ�1�C���g��� ��ߘ���P���t�	� ��?���c�u��� (����^������� $�M���q� �����6� ��Z�����%��I [���2��~��VISBCK��|��ų*.VD�|*� FR:\�V� Visi�on VD fileVd���� ���	/./�R/� v/�//�/;/�/_/q/ ?�/*?<?�/`?�/�? ?�?�?I?�?m?OO �?8O�?\O�?�?�O!O �O�O�O�O{O_�O!_ F_�Oj_�O�_�_/_�_�S_�_w_�_o~�MR_GRP 1=���LeC4  ;B�`	 ��lo�~li`۬B���D��fn�ӺMT� �?�� ����e`i `a�o�khb�h�o�d�cic.N�d�4L7>K�4��M��HC�E��|�i`�@
�B����A�h?
�7�BX=�9�h�l}A�b�A����A��A�I_�A辊�p�l}F@ �qhq�y�~�g�fF6�D��MqD�� BT��@���l}�?pD��6����l���5���5��|��~e9��B�yA��bA�	m�zsA�-G*eA����z󏶈������A�܏e�P���t�  �@߬�?R�Z�?AZ}@�rS �����Ο��+�� O�:�_���p�����veBH` �x����a;�ީ����'�d
��Z��WZ�!/�FX�
�A@����@�3w3@����\��[���ѿ�z��񿋯 �*��N�9�r�]ϖ����<�G�=��<�m]<��+=~�m<c�^��8eN7���7ѷ7��x7;��51�@��	ߤ��?߾d2^`UYb`�b`��������F�`Үb` b`:��0�����C�^o �߂o�o�߸o��o��  ]�(߁�l����� ��������#��G�2� k�V�{����������� ����1 �� -�)����� ��0T?xc �������/ ')�'/M/_/q/8��/ �//�/�/�/�/?#? 
?G?2?k?V?�?z?�? �?�?�?�?O�?1OO UO@ORO�OvO�O�O�O �O��_��J����`_ *�_N�_�O�_�_�_ �_oo'oMo8oqo\o �o�o�o�o�o�o�o �o7"[Fjh �x�t��!�� E�0�B�{�f�����Ï ���ҏ����A�,� e�,/���������/� J����=�$�a�H� Z���������߯ʯ� ��9�$�]�H���l� ����ɿ��ƿ���#� �O�OV� _z�D_V_�� z_�Ϟ_���
�C� .�g�Rߋ�vߛ��߬� ����	���-��Q�<� N��r������� ���)��M�8�q�\� �������������� ��7"[Fk�| �|����֟3 �WBg�t�� ���/�///S/ >/w/b/�/�/�/�/�/ �/�/??=?(?:?s? :�LϦ?p��?�Ϧ� O ��$O��T?]OHOZO�O ~O�O�O�O�O�O�O_ 5_ _Y_D_}_h_�_�_ �_�_�_�_�_o��@o 
�go*owo�o�o�o�o �o�o	�o-*c N�r����� ��)�;�M���� �����ˏݏď�� %��I�4�F��j��� ��ǟ���֟��!�� E�0�i�T���x���ï �?�?��O��?OO �t�>O������ѿ�� ο��+��O�:�s� ^σϩϔ��ϸ����� � �9�$�6�o�6o�� Zo��R���������� 5� �Y�D�}�h��� �����������
�C� U��y�����d����� :�����+Q8 u`������ �;&_Jo ������// گ4/��x�j/4��/X� n/|��/��/�/!?? E?0?B?{?f?�?�?�? �?�?�?�?OOAO,O eOPO�OtO�O�O���O �O_�O+__O_:___ �_p_�_�_�_�_�_�_ o ooKo6oooZo�o Z��o�o�o�o��xo 
G2kR��� ������1�� .�g�R���v�����ӏ ���	��-��Q�/ */��N/��r/�/ޟ�/ ��/)�D�M�8�q�\� �����������گ� ��7�"�[�F�k���|� ����ٿĿ���O�O�O ��W�B�{�fϟϊ��� ����������A�,� e�P߉�t߆߿ߪ��� �o��+�=�a��� ��p���������� � �9�$�]�H���l� ��������������# G2W}h�p���$FNO �������
F0� ��  #�1 D|��� RM_CHK�TYP  � �\q�� �� ��{OM� _MIN� �m����  �X� SSB_C�FG >� ~�Jl��Aj|�TP_D�EF_OW  �m���IRCO�M� ��$GENOVRD_DOs����THR� d�d�_EN�B� �RAV�C_GRP 1?3� X�e/� �/�/�/�/�/�/�/�/ ? ?=?$?6?s?Z?�? ~?�?�?�?�?�?O'O OKO2OoO�OhO�O�O��O�O�O�O�ROUr? E� q�������8�?#�O__K_m_o_�?�  D3���_�E�_q�@A��\B�����R��>Y_6 SMT<#FC-�Ufoxo|�o�HOSTC,s1GY?��_k 	�h�k�o2�f�oyeC Ugy�z1�������p	ano?nymous�5� G�Y�k�w��o�o�o�� ����*�<�� `�r�������ˏ	�� ���&�8������� �������ȯگ��� M��4�F�X�j����� ݟ��Ŀֿ���I�[� m�ρ�fϵ��ϜϮ� ����}�����,�O� Pߟ�t߆ߘߪ߼�� �/�A�C�(�w�L�^� p����ϸ������� ���a�6�H�Z�l�~� ����������9�  2DV��z�� ����#��
. @������������ ���//g</N/ `/r/�/����/�/ �/?Qcu��/[? ��?�?�?�?�?)/�? O"O4OFOi?�/�/�O�O�O�O9m�aENT� 1H[ P!\^O_  `_ ?_._c_&_�_J_�_n_ �_�_�_o�_)o�_Mo oqo4o�oXojo�o�o �o�o�o7�om 0�T�x��� ��3��W��{�>� ��b���Տ������� ��A��e�(�:���^�𿟂�㟦�QUICC0�̟ޟ?��A1@��.����2���l�~�߯!ROU�TER௼�ί/�!?PCJOG0���!192.168.0.10	���GNAME !��J!ROBOT����NS_CFG �1G�I ��Auto-s�tarted/4FTP:?�Q?SO Bχ?f�xϊϜϮ��? �������+�߿�P� b�t߆ߘ�6��� ��(�J� �1�C�U�g� 6ߋ���������x� 	��-�?�Q�c� ?2? D?��������� )��M_q���� :���%t� ����m������ ����!/3/E/W/ z{//�/�/�/�/�/ 6HZ ?n/S?�w? �?�?�?�?�/�?�?O O<?=O�?aOsO�O�O �O�/
??.?0O_d? 9_K_]_o_�_PO�_�_ �_�_�O�_�_#o5oGo Yoko�O�O�O�O�_�o &_�o1Cog y����oT�� 	��-�|o�o�o�o� ���o��Ϗ���� )�;�M�_�q������๟˟ݟ�ÿT_ERR I������PDUSIZ  ��^���$�>~=�WRD ?޵�w��  guest+�}���࡯��ůׯ��SCD�_GROUP 2]J� �`�51��!��L_����  ��!�	 �i-	�E����Q�E EATSWILIBk�+���ST 4��@��1��L�F�RS:аTTP_AUTH 1K��<!iPendCan�������!KAREL:q*���	�KC��.�@��VISI?ON SET���u���!�ϣ������ ��	��P�'�9߆�]��o޽�CTRL �L��؃�
���FFF9E3���u���DEFA�ULT��FA�NUC Web �Server��
 ��e�w���j�|���������WR_CONFIG MY�X����I�DL_CPU_P5C���B�x�6�w�BH�MIN'���;�GNR_IO��K���"��NPT_SIM_DOl��v�TPMODN�TOLl� ��_P�RTY��6��OL_NK 1N�ذ �� 2DVh��_MASTEk�s��w�OñO_CFG���	UO����C�YCLE���_?ASG 1O��ձ
 j+=Oa s�������p//r�NUMJ�� �J�� IPCH��x��RTRY_�CN�n� ��SC?RN_UPDJ�����$� �� �P��A��/���$J�23_DSP_E�N~��p�� OB�PROC�#���	J�OG�1Q� �@��d8�?р +S? /?)3PO�SRE?y�KANJI_� Kl��3��#R�����5�?�5CL_LF�;"^/�0�EYLOGGINʦ q��K1$���$LANGUAGgE X�6��Y vA�LG�"S��V������x��i�j�@<𬄐'0u8������MC:�\RSCH\00�\��S@N_DISP T�t�w�K��I��LOC��-�D�zU�=#�J�8@B?OOK U	L0���d���d�d��PX Y�_�_�_�_�_ nm1h%i��	kU�Y�r�UhozoLRG_B�UFF 1V��|o2s��o�R���o q��o�o#,YP b�����������(�U��D/0D�CS Xu] =���"lao����ˏ�ݏ�3n�IO 1Y	 �/,����,�<�N�`�t����� ����̟ޟ���&� 8�L�\�n����������ȯܯ�Ee�TM  [d�(�:�L� ^�p���������ʿܿ � ��$�6�H�Z�l��~ϐϢύd�SEVt� ]�TYP��$���)߄m�1R�SK�!O�c�"FL 31Z�� ����߀����������	�:�T�P5@���A]NGNAM�$�E��k�7UPS PGI|%�1��%x�_LOAD�0G %Z%0_MOV�e����MAXUALRM ;'�I(��~���#� QV�#a��CQ[x�@8��n��"�1060\	 �F�	�Ϣ��� ���������� D '9ze���� ����R= va������ ��*//N/9/r/�/ g/�/�/�/�/�/?�/ &??J?\???�?k?�? �?�?�?�?�?�?"O4O OXOCO|O_OqO�O�O �O�O�O_�O0__T_ 7_I_�_u_�_�_�_�_��_o�_,o��D_L?DXDISAc����MEMO_AP�]�E ?��
 �5i�o�o�o�o��o�o�o��ISCw 1]�� �o Td��\no�� �������I� 4�m��f���$����� ����!��E�ƏT� f�:�����ß����� z��ܟA�,�e�w�^� �����~������  �=���L�^�2����� ����߿�r� �Կ9��$�]�o�(t_MST�R ^�͂�SC/D 1_xm�W��� S�������=�(�:� s�^ߗ߂߻ߦ����� ��� �9�$�]�H�� l������������ #��G�2�W�}�h��� ������������
 C.gR�v�� ���	�-Q <u`r���� ��//'/M/8/q/�\/�/�/�/�/�/s�MKCFG `����/��LTARMu_2a��2� �#\`Y>G`M�ETPUT`�"�����NDSP_CMNTs506�5��' b���>�"1��?�4�5POSCFz�7�>PRPM�?��8PSTOL 1�c2}4@p<#�
aA�!aEqOG]OO �O�O�O�O�O_�O�O A_#_5_w_Y_k_�_�_�_�_�Q�1SING_CHK  +O�$MODAQ73d�
?�7:eDEV �	��	MC:>MlHSIZEs0����eTASK �%��%$1234?56789 �o�e�gTRIG 1en�� l��%��?   A$�Üf�YP�a,u��cE�M_INF 1f�>7 `�)AT&FV0�E0N�})�qE�0V1&A3&B�1&D2&S0&�C1S0=�})GATZ�� �H� E��q9m��xAu��� X�������� �� ����v�)���я ��П�������*�� N�����7�I�[�̯ ן���9�&���\� ���g�����i�ڿ�� ����ï4��XϏ�i� ��A���m�������� ��ѿB����ϊߜ� O������ߟߩ���� >�%�b�t�'ߘ�K�]� o߁�����(�_�L� ��p�+����������.�ONITOR�0G� ?ak   	?EXEC1�#U2345T�`789�#��xxx *x6xBxNx@Zxfxrx2U2�2�2�2�U2�2�2�2�U2�33�3�aR_GRP_SOV 1g�y�a(�Q�?i=�?�vq���	@M���
�y<�Hm�a_Di�n�!P�L_NAME �!�5
 �!D�efault P�ersonali�ty (from� FD) �$RR�2� 1h)de�X)dh�
!�1X d�/d/v/�/�/�/ �/�/�/�/??*?<? N?`?r?�?�?�?�?�?�82S/�?O O2ODO@VOhOzO�O�Ob<�? �O�O�O�O_"_4_F_�X_j_|_�_LhR� �1m)9`\b0� �_pb�Q �@D�  �Q?���S�Q?`�QaAI?�Ez  a@o�g;�	l�R	 O0`4b@4c�.a�P�Jd�Jd�K�i�K�J����J��J�4�J~��j0Ea�o-a�@��o�l�[`@�z�b�f�@�S��a�Q�o��c�=�N��
������T;?f�
���m[`��*  �p  ��$p> p�$p���o?��?�����	��o�Bntr�Q�s�kse�}�l�p��  �pu`j7  #p��vks��� 	'� �� �I� �  ���}�:�È6�È=����N��b@�^�d��n�Q���{�RȒx���nN. ��  �'���a�`@a��@�t�@p@hp�n[`CpC0��f0�+pB/pC3}��P�@%�Ea�  oo�$|m����gA%���. ���z!�`�P���QDe����˟��(��m��� �t O�� ru �4 �R�c��sO� :	e�a�P~�` �?�ffd��!�����7� ���گ쬛af��>搠���iP�P;�e��S�Ea4f�u�>L�X��s�b<	�I<�g�<#�
<�2��<D��<���
vo��¯�S���S.���?fff�?u�?&찗d@T����?�`?Uȩ?X�� ��Z���T:z�TB��W a�з*dů�ρϺϥ� �������&�8�#�\�h�+�F. Kߘ�G߀��3���Wɯ���G?�@ G���� X�C�|�g�y����� ����jZ���ￏQ� ���ߙ�����3��� ����/A��t�_������� ����d���@+Fp�IP�t�e�%���[`B�0� ���<ze�cb�!@I�
�M`�B@��@`��9@y��?��h� �@�3��[N��N�N��E��<�/�:/L �>��ڟ��A�p�C��F@�S�b/�X������@��t��%�h���`/qG��G�knF&�F׿�pE,8{�/ �F�ZG����F�nE��DE,ڏ�/� ����G��F7���F��ED��.��C?.?g?R?d? �?�?�?�?�?�?	O�? O?O*OcONO�OrO�O �O�O�O�O_�O)__ M_8_q_\_�_�_�_�_ �_�_�_o�_7o"o4o moXo�o|o�o�o�o�o �o�o3WB{ f������� ��A�,�Q�w�b��� �������Ώ��� =�(�a�L���p�����=(r!3�ji��r����ꕢ�3Ա�xڟ�u�4 ���<�u�P�2�D��&�jb^�p�1w?����������ʯ���ܯ� �s�P^�PD�c�`�m���@y�\������Ӱ�¿ Կ�����.�G� ���}ϳϡ���홍�@U�_�J���$�y.� @�v�d�z߈ߚ�x�4� �������� ��D�.��2� �$[�G�D[�^�B���B��CH� ^����u��@��������p�h�M�_�q�����������^�^�Y�m�2��
 ���� #5GYk}�������h*�� ���>�x}��$�MSKCFMAP�  ��� ����m�N"�ONREL  �6�9_�"EX_CFENBk
7�]�FNC�}JOGOVLIMk�duyd"KEY�k�"RUN���"SFSPDTYU��v_�SIGNk}T1�MOT�z"_�CE_GRP 1-n��9\���/ ���/�/4��/?�/2? �/'?h??�?C?�?�? y?�?�?�?O�?@ORO 	OvO-OoO�OcO�O�O �O_�O*_<_#_`_-��"TCOM_CF/G 1o/���_��_�_
|Q_ARC�_�6��UAP�_CPL�_�NO�CHECK ?/ 5�;h9o Ko]ooo�o�o�o�o�o �o�o�o#5GT�NO_WAIT_�LF'5y"NT�Q�p/���q_ER�R�!2q/_�� AR_���"�x:�L�dT_MO�s}r�}, ��.P_|��_�PARAM�rs/�������MW��� =e�345678901.� @�R�)�q���_������˟����ݛLW��3�E�؏i�cUM_?RSPACE,��������$ODRD�SP�SI&�OFF�SET_CART�oݨDIS�ݢPEN_FILE��I!�Q�v�POPTI�ON_IO���PWORK t�'� T�|�/�^��F�U��Z���	 ��m���C�����R�G_DSBL  ���v���ޡR�IENTTOj���C���8=#��?�UT_SIM_EDJ�6	��Và?LCT u�}�\��Q��W�_PEX9E���RAT���� ���UP )ve���������X��*�8��$��2�#�h)deX)dh}�O�X dY� ߑߣߵ��������� �!�3�E�W�i�{��@�����������2n� �)�;�M�_�q���������<����� +=Oas��ЩX��� O��1m(���(�.��g��"0 ��дu�  @D� M �?��?р�H�D4  EzxZ3;�	l?	 0ӀSQ@SM� �i�i� �H)!H,��H8�Hm��G�	{G�81��6�MV���� �C�)���)�����Ճ�*  ��p  � > �  ��/$"��,��B,�Btr߰«�H�¼�/���/�"`�# �,0 �� _�  � ߽poj   ��&�X�?MU	'� �� 12I� ��  ���-=����U?g;/�@}?�0~.ѱ�?;Ѳ1���H[N �?Aa'M�D�> C)�	f)�" B& �"O4Bx+�:�Q�@D1~�oo$�����JWA�D0�J@�A:  �1�E&?�O�O#_�_G_2]�� ��t O� �ru �4 ���R�Uɳ� :��%S�р� �?�ff��@[�_�_BV_{�o~��18р�"o0j>�P�Q6YP�рZo�WrAdS�%��>Lw0�#�<	�I<g�<5��<2��<D��<�ל���_�j��ѳMb�@?ff�f?�0?&p:T@�T�q?�`�?Uȩ?X� -q�iyBq5Ya ��gI�_��� ���!��E�W�B� {���d�����ՏLn�pΏ/�ʈG�@ G��U�ȏy�d��� ����ӟ������� yB=� ��?p���/� ���߯R���'�9� �oN�`�����~�����ۿƿ�B�ĮD��e�ֿ;�ҿ_�J�?Ƀ�h�oϨϓϸ��D4��b!�_@����� ߧ��Ŀ����%�@�I�)�M`B@���@`�9@y��?�h	�� �@�3�[�N��N�N�E?��<�/Y�k���>��ڟ�A��p�C�F@�S���pX������@�t�?�%�h��߉!�G��Gkn�F&�Fצp�E,8{�� F��ZG���F��nE�DE�,ڏ��ૐ��G��F7��F��ED��Mf ��b�M��q���� �������(��8�^� I���m����������� ����$H3lW �{����� �2VAS�w ������/./ /R/=/v/a/�/�/�/ �/�/�/�/??<?'? `?K?p?�?�?�?�?�? �?O�?&OO#O\OGO@�OkO�O�O�O�N(]��3�ji�O�a��<	U�E3Ա��O_<q4 ��%_7_<q��P�Q_c_ER�jb}_�_1w������]�Y�_�_�o�_1ol��P�bPcn~���o�O�o{_�o�oY�`��o�o, /;M#�f0o� ����Y�et�~�i#�1�C�yM�_��� ��������{bS�Ԏ�@�	�?�-�c�Mj2��;�$�VG�z}��B����B��CH �}�9�֟�����0�B���wl�~���P����Ư�T�퀑�\��qQ��U
 ί�0�B�T�f� x���������ҿ����χ��� ��]{x�}��$PAR�AM_MENU �?Յ��  DE�FPULSE��	WAITTMO{UTl�RCV�� SHELL�_WRK.$CU�R_STYLj����OPT����P�TB����C��R_DECSNw�Te'� !�3�E�n�i�{ߍ߶� ������������F��A�USE_PRO/G %P�%B��.V�CCR��UeX����_HOST �!P�!�����T t`���������4�>��_TIME�� ��T�  A�GDE�BUG��P�V�GI�NP_FLMSK�]���TR����PG�A�� |�[���CyH����TYPEM�Y�A�;�Qzu ������
 )RM_q�� �����/*/%/ 7/I/r/m//�/�/�/��/�/?��WORD� ?	��	RyS��CPNS�E���>2JO���B�TE���TRAC�ECTL�PՅ�Z� {`* +�a`{`�>q6D/T QxՅ�0�0�D�� #����0���2&�4'z��Sc{a��0��B�� �5�0�2�0B�0B�0P��2��2�4�4U	�4�4�4�4E�4�4 ��2�4U�4�4�4�4U�4�4�4�4��2�4�4���2!�4"�4�?�8DOVO hOzO�O�O�O�O�O�O�O
Z%�9O.O@O2_ D_V_h_z_�_�_�_�_ �_�_�_
oo.o@oRo dovo�o�o�o�o�o�o _V!3EWi {��������5�( �)�"�4� F�X�j�|�������ď֏��1u�*� <�N�`�r��������� ̯ޯ���&�8�J� \�n���������ȿڿ ����"�4�F�X�j� |ώϠϲ��������� ��0�B�T�f�xߊ� �߮����������� ,�>�P�b�t���� ����������(�:� L�^�p����������� ���� $6u� bt������ �(:L^p ������� / /$/6/H/Z/l/~/�/ �/�/�/�/�/�/? ? 2?D?V?h?z?�?�?�? �?�?�?�?
OO.O@O ROdOvO�O�O�O�O�O �O�O__*_<_N_`_ r_�_�_�_�_�_�_�_ oo&o8oJo\ono�o V�o�o�o�o�o�o "4FXj|�� �������0� B�T�f�x��������� ҏ�����,�>�P� b�t���������Ο�� ���(�:�L�^�p� ��������ʯܯ� � �$�6�H�Z�l�~��� ����ƿؿ���� � 2�D�V�h�zόϞϰ�������$PGTR�ACELEN  ���  ��������_U�P y���2�������_CFG z�S������<��� <�Z�l�<�$��DEFSPD e{/��a������IN'�TRL �|/���8Lԃ�I�PE_CONFI�+�}��t�<�x�LID(��~/��GRP s1���������@�
=�[����A?C�C
��XC)��B�Y�r������dL��z������� 	� r�N��Ҩ�� #´����B�����������A���> �6>7�D_�������� ='�=)��������� 	B-��Q�Mx���  Dz����
��&L 7p[���� ��/�6/!/Z/���
V7.10b�eta1<�� �B=q�"`ff�@��">���ާ!=��͏!A>{ff�!@�ff�"��\)�"D��?�  �!@�!� �!Ap�#W��h/??*?<?K;�w����O/�?K/�?�?�?�? O�?O>O)ObOMO�O qO�O�O�O�O�O_�O (__L_7_p_[_m_�_ �_�_��_ o�_$oo !oZoEo~oio�o�o�o �o�o�o�o DQy<{/�#F@ {yw} �y{ջy�-��� ���/�Z?l?~?w��� t�����я������� ��O�:�s�^����� ����ߟ�ܟ� �9� $�]�H���l�~����_ ۯ�����5� �2� k�V���z�����׿¿ �����1�\n�j� |϶�������	� 4�F�X�j�c�χߙ� �߽ߨ��������)� �&�_�J��n��� ��������%��I� 4�m�X�����ί���� ������!E0B {f������ H�Zό�Vh�� �ϊ����� �2� D�V�O/�s/^/�/�/ �/�/�/�/�/? ?9? $?6?o?Z?�?~?�?�? �?�?�?O�?5O OYO DO}O�O���O�OtO�O �O_�O1__U_@_R_ �_v_�_�_�_�_�_" 4FxBo|��� �o��o�o//0/B/ ;�__J�n�� �����%��I� 4�F��j�����Ǐ�� �֏�!��E�0�i� �O^���N�ß՟���� ���A�,�e�P�b� ���������o o2o To.�hozo�o�����o ��Ϳ�o
گ'�֯ K�6�o�Zϓ�~Ϸ��� ���������5� �Y� D�Vߏ�z߳ߞ����� �����1��Uy� ��:���������	� ��-��Q�<�u�`�r� ���������� T�f�x�n����� �������7" [Fj���� ���!//E/0/i/ T/f/�/�/�/�/�/�/ ?�//?A?l�e?w?&? �?�?�?�?�?�?�?O O=O(OaOLO�OpO�O �O����*�O_@R�dZ_l_��$PL�ID_KNOW_�M  ����A�TSV ����P�[?�_�_o�O�&oo#o\o�B��SM_GRP 1��Z�� dI`�o�o$Cf�d����D��TPbj �oLk�f�o"~�U�o> n2T�~� ����7�4��� p�D���R���ʏ���� ������6�
�T��*�X�����QMR�c��m1T�EGQK? GR� �(�#���[��/�A� S������������$� ���W��+�=�O��� ��������� ����S�Ͻ�ST�a1 �1������P0� @����E�� ����������M�0� B�T�fߧߊߜ����� ������7��,�m���2�����A�<��z�3�������A4���������5)�;�M�_���6x���������7�����������8(:L��MA/D  ���� ���PARNUM � ��Ko���S+CH�
 �
�8�S+UPD���xaq{��_CMPa_�`� <Pz '�U~�ER_CHK�����Z���RqS���_�Q_MO� ��%_��_REWS_G����� � �v/{/�/�/�/�/�/ �/�/*??N?A?r?e?w?J'��W,g/�?L% ��?�?�?N#(��?O ON#w�4OSOXON#�� sO�O�ON# �O�O�O�N#d �O__N"V �1��Uua�@cX���Pp�P$@cW�،P��P@@cV���P�"THR_�INR���pbA%dޠVMASS�_ Z��WMN�_�SMON�_QUEUE Q��e��`Ȩ`�N�U�N�V�2`�END4a6/NiEX1E]oNeWBE\`>o>/cOPTIO;g?+�2`PROGRAM7 %j%1`O_��0bTASK_I���nOCFG �o�9pDATuAɓ�B{@ev2w������z� �+�=�O��s�����x����nzINFOɓ��}�!dr��!�3� E�W�i�{�������ß ՟�����/�A�S��e�w�҇ބ��| ��98q�DIT �Bׯj~WERF�L~hwS~�RGAD�J �ƪA� � ,�?E�8��Q�I�ORITY�W��>�MPDSP�a��j�U�WvT�OG��_TG���Rj���TOE�P1�ƫ� (!AF�PE�5 ���!tc�p��%�!ud|�?�!icm<��Q_��XY_<q��Ƭ�Oq)� *0������Op����� �������<�#�5�r� Yߖ�}ߺ��߳�������&�*�PORTT�a�OpA%��_CARTREP�~`Ʈ��SKSTA��X!*SSAV`��ƪ	2500H809u�T毙䕣U�ƫ�����`�X#�$�6�m�URGeEU`B��A)WFP�#DO�V�2�W�q��?Q�WRUP_DELAY �Ư>e�R_HOT�hwR�%z����R_NORMAL�n��6SEMI:y�_QSKIP���X%;�x 	��� �����X%- ;%[mE�� �����!//E/ W/i///y/�/�/�/�/ �/�/?�/?A?S?e? +?�?w?�?�?�?�?�?�O�?+O=OOO1U�$�RBTIF��NaR�CVTM������m@DCR�����A;��BI��Y@�Y?���ۧ�=�|���}`��uH��'_S<	�I�<g�<#�
�<2��<D��<��
+__{_�_ )`���_�_�_�_�_ o o$o6oHoZolo~oi_ �o�o�o�o�o�o�o  DV�_z��� ����
��.�@� R�=v�a��������� ��׏�*�mN�`� r���������̟ޟ� ����8�J�5�n�Y� ��}���ȯ�����A� "�4�F�X�j�|����� ��Ŀֿ�ӯ���0� B�-�f�Qϊ�m���� �������,�>�P� b�t߆ߘߪ߼ߧ��� �����(�:�%�^�A� ����ϸ������� � �$�6�H�Z�l�~��� {������������  2Vh���� ����
.@ R=O�s��� ��/�*/</`/ r/�/�/�/�/�/�/�/�??&?28�AGN_�ATC 1��K� AT&F�V0E02;A�TDP/6/9/�2/9p8ATA�2>,AT%G1%B960k9_+++�?,�1�_,�AIO_T?YPE  EC�/4?REFPO�S1 1� K 'x�O[H/O /�O�MNO`O�O�O�O _�OC_�Og__d_�_^+K2 1� KLO�N_�_o�_*o�_5A3 1��_�_�_ o�o��o�o@oS4 1� Woio{o�o3W�oS5 1��o�o�J���jS6 1�����]�H�|���S7 1���(�:�t��ݏ���S8 1�����Ϗ	����r���)�SMAS�K 1� O  
8���ɗXNO�?����1.�8�1AMOT�E  �.DN�_CFG �U���5��0BPL_RANG�Q�K!Y�POWER� �Q5 a�S�M_DRYPRG %�%R���ȥTART �����UME_PRO�ׯ�d�.D_EXE�C_ENB  <�5]�GSPD=��8��Y3��TDB����sRMÿ��MT_ѐ�T��S�D0OBO�T_NAME ��S�;9OB_�ORD_NUM �?��A�H80�0I$�	/��s	�\���{�� ��e��7	@�}�D|��D0�PC_TIMEO�UT�� xD0S2�32n�1�Q; �LTEACH PENDAN���j�5��=Q�x0�Maintena�nce Cons�K"-��"+�t4KOCL/C�}�6���|� No Use�=[߹�Fώ��NPO�ќ�5��_���CH_�L@��U���	�J��MAVAIL�`���+��]�I�SPACE1 2�=L ����p���扢J@����8�?��� ��� V�w�N����������� ����4�&G
l� }d	Q5U1������� ��`4&G
l�}d�#��2�� ������2A/�b/%/w/�//�/�3 ����	/�/-/O/ ^??B?�?�?�?�?�4�/�/??&?�?J? l?{O�O_O�O�O�O�O�5�?OO1OCO�O gO�O�_�_|_�_�_�_o�6_*_<_N_`_ o�_�_�o�o�o�o�o!�75oGoYoko }o+�o�o����)��>��8Rdv ��H�����ӏ�%�F�-�[��G ��� R�;�
�� ����ԟ� ��
��.�@����c�@��p���8�¯=�dؠ ��ϟ���!�3�E�W� i�_�q������x�� կ��'�9�K�]�o� ��w��ϛ���Ͽѿ� ���5�G�Y�k�}ߏ߀�ߗ��߻������; `S� @��8�@��F�"�*ل��� ���߇������ ,����V�h�2�<�N� ������������. L4v�R\n�����
f�7��_MODE  ���MS ���&����Ïb���*	�&/�$CWO�RK_AD]�{�x�!R  ����t +/^ _INOTVAL]���h�R_OPTION��& h�$SCAN_TIM\�.�h�!R ��(�30(�L8�E�����!��3��1�/@>.?V���S22�4D11d�8�1�1"3��@���?�?�?����IP����@���JO\OnOE@D���O�O�O�O�O �O__(_:_L_O���4X_�_�_���8�1��;�o豔 1��pc]�t��Di�1��  � lS2��1 5 17oIo[omoo�o �o�o�o�o�o�o! 3EWi{��� �wc���	��-� ?�Q�c�u��������� Ϗ����)�;�M� _���`[����ğ֟ �����0�B�T�f� x���������ү���p��$�7�  0� �� om��������ǿ ٿ����!�3�E�W� i�{ύϟϱ������� v���/�A�S�e�w� �ߛ߭߿�������� �+�=�O�a�s��� ��ߖ����� ��$� 6�H�Z�l�~������� �������� 2DVP�\�  �A�� �����% 7I[m��������/ � /C(/N/`/r/�/�/��/�/�/�/�/?F�;/?B?F�x1� ;?w=	12�345678{���l�@��P�?�?�?�?�?O 9/2ODOVOhOzO�O�O �O�O�O�O-/
__._ @_R_d_v_�_�_�_�_ �_�O�_oo*o<oNo `oro�o�o�o�o�_�o �o&8J\n ���o����� �"�4�F�X�j�|�� ����ď֏����� 0�B�T�f��������� ��ҟ�����,�>� m�b�t���������ί@����(��6y I�[�@�`���������Cz  Bp*_   ���254�F��$SCR_G�RP 1�(�e�@(�l�}�0@ `1� [1s	 )� 3�C�<�t�vrY�8�P�}�kϤ�����95C����-u���ȡ���LR �Mate 2007iC �190�1�~�0LR2C �3P�=OÆ�D�
f��1u�2�U7��`1��Dv��@�u���	t�@��������$�^0�2���_2T�gϡ� ���o�F�D�f?��s������￶ht ,Z��r�B�˰ƐP�N�g�N�Aܰv� # @DЎ�N�@����G  ?� ��J�H˰���y�N�F@ F�`������A ,Qwb���n� N�������B��_J�n �����/�%/ /I/��E+:3��6?|?��5��
�/�/�#��@=��"�/pǢ�� 3B�07�59�0@7���EL_D�EFAULT  �I����� ^1MIPOWERFL  V�xv5]2�0WFDOk6� v5 �ERVE�NT 1����O�t3C�L!D?UM_EIP?�8��j!AF_I�NEj0O�$!FIT�?=NOaO!Q�ΆO �PO�O!�RPC_MAINĮO�H��O�O�CVI�S�O�I��OE_!�TP8PPU<_�9d�4_�_!
PMON?_PROXY�_�6Ae�_�_XR�_�=f�_�)o!RDM_S�RV*o�9gouo!#RR8�o�4hdo�oK!
�@M�_�<i�o�!RLSYN�C4y8�oY!�ROS�?�|�4 H�tO�8c��� ��;��_�&���J� ��n������ȏڏ 7�I��m�4���X�����7ICE_KL �?%�; (%SVCPRG1�� ���!��3*�/�"�4R�W��5z��"�6�����7ʯϯ��C��5�9�� oG����o��� ���D����l��� ���񑼯7���_� �����4����]� ����������'�� տO����w��%ϟ� �M����u������ ����?�A��Ͽ�ђ �؟ꐊ���ɱ���� ����?�*�c�N��� �������������� );_J�n� �����% I4mX�|�� ���/�3//W/ i/T/�/x/�/�/�/�/��/�/?/??S?Ś_�DEV �9��MC:[8��im4OUT_R�f1~6i8REC 1q���f0�0 f0_ 	 f0�2  
f0�4�1���3OMK�1�4=A�%O^OAA��
 �Z�6 s;B �3AAqE=�=A���2WG��1f0)f0{f0U��Of2B0����	�/Q0�O_�5�媂@��@r�H�;@��  x�0}@ZU@��O f0�f4J�1af0�V_�2X0U��@�f0?�@�~_��__��2\�0���0��0�@�����_ f0�f0�1=Jf0[f0�o�2T0U��@�f0*�@u*o,co�_�ÆLH�0�0���R �  ��RobmU�f0z�f0�o�2�Q��@ъf06�@z�ovo~QK�L=A�1(f0tf0�f0�_c�f4e�=ѭZZ f0k0�*�0Cf0f0q��"~N�LiI�1�2��f2Pf0>jI��zD�f0f0o.�g���UφL"f0i�0bf0���0��0V�b��f0f0/f0|~ �0��E0��@��f0$�@Y�^�p����B�L*�A�0=�QpɀS��b�ʈ�f0�_^�f2C0��@���A0����&���2\�AM��Up���A��p�<~��O���b��$2�k�ҟ�2\i&f0}��0�0�Wf0�Z��b�f0Jf0R~�[���F��@	ݒq0"ޯ�*�a @��Z�H�~�l��� ����ؿ������2�  �V�D�zό�nϰϞ� ����������.��>� d�R߈�v߬ߚ����� �����*��:�`�N� ��f�x�������� ��&�8��\�J�l�n� �������������� 4"XFh�p� �����0B $fT�x���<��5V 1��<���`!	O�2 W��P���a?�_TYPE�?k2H�ELL_CFG ��z:f2/ 8HL�/<7RSա�/ �/�/"??F?1?j?U? �?y?�?�?�?�?�?O��?0OBOQK��p�!%QOO�O%��x�q`�qQ��M�q�p�$��gBQ�d�O�O�&HKw 1��+ �O E_@_R_d_�_�_�_�_ �_�_�_�_oo*o<o�eo`oro�oa&�#OM�M ��/�o�"F?TOV_ENM�t"�!}*OW_REG�_UI�o�"IMW�AIT�b���G${O�UTv$&yTI�Mu��`VA�L5's_UNIT��c�v})MON_ALIAS ?e�i? ( he!�  ��$�6�%��c�u� ����D���Ϗ��� ��)�;�M�_�q���� ����˟ݟ����%� 7��H�m������N� ǯٯ������3�E� W�i�{�&�����ÿտ 習���/�A��e� wωϛϭ�X������� ����=�O�a�s߅� 0ߩ߻����ߊ���� '�9�K���o���� ��b��������#��� G�Y�k�}���:����� ������1CU  y����l� �	-�Qcu �2������ /)/;/M/_/
/�/�/ �/�/�/v/�/??%? 7?�/[?m??�?<?�? �?�?�?�?�?!O3OEO WOiOO�O�O�O�O�O �O�O__/_�O@_e_ w_�_�_F_�_�_�_�_ o�_+o=oOoaosoo �o�o�o�o�o�o '9�o]o����P������s��$SMON_DE�FPRO ����:�� *SYST�EM*  �l��*�RECALL� ?}:� ( ��}Ecopy �md:cal_d�v_xy.tp �virt:\ou�tput\��ov�er =>330�30144:694973�Џ⏻pc}9z�����ls~� ������E�W��y��� ������ҟ���	�� -��P�b�u�������=�ί��;z�fr�s:orderf�il.dat��t�mpback\=�>laptop-�3jv248ms:��48 ��G�Y���2z�b:*.* �!�3�-�f�п���6x��:\����������B�T��7��a���+�2������8����z�����D�V�
�Cz�z�����;� >����������*��� G�Y�l�~�4��� ������� ϲ�C�U� h�z�����6������l��ς�ptcp.pcߴس�DV�5�� _1��2 ��hz�2�� �FX����_� &8���Az� ��&�+�P/b/u �,�3/�/�/�� �+/�/B?T?�/��� �ﯴ6?�?�?l�~�? ��?EOWO����� � 2O�O�Oh/z��O�O�� �OG_Y_�/�/?��0_ �_�_�_x?�?O.O?o Qoco�?o#o,O>o�o �otO__�O�oM_ �O(_:���_ o�o&o�I�[�no�o ��o6�Ǐُ�o�o� "��E�W�j|�� 2�ß՟h_z_�_�_�� A�S�e�x/���6� ǯٯ����"��E� W������2�ÿտ h�z�������A�S�e���$SNPX_A�SG 1�������� �P 0 '%�R[1]@1.Y1fϰ�?�p�%�� �Ͽ� �����6��@� l�Oߐ�s߅��ߩ��� ���� ���V�9�`� ��o���������� ���@�#�5�v�Y��� ������������ <`CU�y� �����&	0 \?�cu��� ��/�/F/)/P/ |/_/�/�/�/�/�/�/ ?�/0??%?f?I?p? �??�?�?�?�?�? O ,OOPO3OEO�OiO�O �O�O�O�O�O_�O _ L_/_p_S_e_�_�_�_ �_�_ o�_�_6oo@o loOo�oso�o�o�o�o �o�o V9` �o������ ��@�#�5�v�Y��� ����Џ��ŏ��� <��`�C�U���y��� ̟���ӟ�&�	�0� \�?���c�u������� �ϯ���F�)�P��|�_�x�PARAM� ����� ��	���P���p�OFT_K�B_CFG  �����״PIN_S_IM  ��̶��/�A�ϰx�RVQSTP_DSB��̲}Ϻ���SR ��	�� & ?CAL_TCŵ�����ԶTOP_�ON_ERR  ������PTN �	���A��RING_P�RM�� ��VD�T_GRP 1�<����  	з�� b�t߆ߘߪ߼����� ���+�(�:�L�^�p� ����������� � �$�6�H�Z�l�~��� ������������  2DV}z��� ����
C@ Rdv����� �	///*/</N/`/ r/�/�/�/�/�/�/�/ ??&?8?J?\?n?�? �?�?�?�?�?�?�?O "O4O[OXOjO|O�O�O �O�O�O�O�O!__0_ B_T_f_x_�_�_�_�_ �_�_�_oo,o>oPo boto�o�o�o�o�o�o �o(:Lsp ������� ���9�6�׳VPRG�_COUNT�q����d�ENB/��_�M��鴖�_UP�D 1�	�8  
M�������-� (�:�L�u�p������� ��ʟܟ� ��$�M� H�Z�l���������ݯ د���%� �2�D�m� h�z�������¿Կ�� ��
��E�@�R�dύ� �ϚϬ���������� �*�<�e�`�r߄߭���ߺ�������\�YS�DEBUGn�Ӏ�� �d��"�SP_PwASSn�B?4�LOG �΅��� ���
� � ��� �
MC�:\`��a�_MPACf�΅����ҁ���� ҁ��SAV ��i���� ����SV�TEM�_TIME 1��΋ (J�;F�0��� ��T1SVGgUNSɀo�'������ASK_OPTIONn�΅�������BCCFG 3�΋O� H�2!`;A�I�r] o������ �8J5nY�} �����/�4/ /X/C/|/g/�/�/ ��,�/�/ ??�/�/ H?3?l?W?�?��?�� �0�?�?�?O�?&OO JO8OZO\OnO�O�O�O �O�O�O_�O _F_4_ j_X_�_|_�_�_�_�_ �_o�X�  o2oPobo to�_�o�o�o�o�o�o �o:(^L� p����� �� $��H�6�X�~�l��� ��Ə���؏����� D�2�h�o������ ԟR�����.��R� d�v�D���������� Я����<�*�`�N� ��r�������޿̿� �&��J�8�Z�\�n� �ϒ���~������"� 4߲�X�F�hߎ�|߲� ���ߤ�������B� 0�R�T�f������ ��������>�,�b� P���t����������� ��(��@Rp� ������ $6ZH~l� ������ // D/2/h/V/x/�/�/�/ �/�/�/
?�/??.? d?R?�?>�?�?�?�? �?r?OO(ONO<OrO �O�OdO�O�O�O�O_ �O__&_\_J_�_n_ �_�_�_�_�_�_�_"o oFo4ojoXozo|o�o �o�o�o�? 0B T�oxf���� �����>�,�b� P�r�t���������Ώ ��(��8�^�L��� p�����ʟ��ڟܟ� $��H��o`�r����� ��2�دƯ����2���P��$TBCS�G_GRP 2���� � �P� 
 ?�  {���w����� տ��ѿ���/�A�T��[��b�d0 ��p�?P�	 HB�HA�L�͌�@�B   C���϶ˀ���ϟ�D����A�(��x���A��T$�9�N�6ff��f�@P�C�ώ�@�f߬��C��ߐ߮ߴޥ��� %��%�D�W�"�4�����j�|�������?Y뙚���	V�3.00s�	lwr2c��	*2��*�O�A� ��ѳ332P�d��� x�J�y�  ������T�JCFG ���l� o������������=K
%�Kq\ ������� �7"[Fj� ������!// E/0/i/T/f/�/�/�/ �/�/�/s���??(? �/[?F?k?�?|?�?�? �?�?�?O!O3O�?WO BO{OfO�O�OP�<��O ��O�O�O0__T_B_ x_f_�_�_�_�_�_�_ �_oo>o,oNoPobo �o�o�o�o�o�o�o :(^L���� ��h� ��$�� H�6�l�Z�|�����Ə ��֏؏� ��D�V� h�z�4�������ҟ ԟ��
�@�.�d�R� ��v��������Я� ��*��:�<�N���r� ����̿���޿ �&� �>�P�b�ϒπϢ� �϶��������4�F� X�j�(ߎ�|߲ߠ��� ��������B�0�f� T��x�������� ���,��P�>�t�b� �������������� &(:p^�� ��t�����6 $ZH~l��� ����/2/ /V/ D/z/�/�/�/j/�/�/ �/�/?.??R?@?v? d?�?�?�?�?�?�?�? OO<O*O`ONOpO�O �O�O�O�O�O_�O_ _&_\_�t_�_�_B_ �_�_�_�_�_"ooFo 4ojo|o�o�o^o�o�o �o�o�o0B�o xf������ ���>�,�b�P��� t���������Ώ�� (��L�:�\���p��� ��ʟ��� ��_�*� �_�l�Z���~����� į�د� �2��� h�V���z���¿Կ� ��
�����.�d�R� ��vϬϚ��Ͼ���� ��*��N�<�r�`߂� �ߖ��ߺ������� 8�&�H�n�\���>� ����x������4�"� X�F�|�j��������� ������
Tf x�D����� �P>tb �������/ /:/(/^/L/n/p/�/ �/�/�/�/ ?�/$?6? ��N?`?r??�?�?�? �?�?�?�? OODOVO hOzO8O�O�O�O�O�O��N  PS �V$_R�$TB�JOP_GRP �2��E�?  ?�W<R�CS�J\��@�0WP�R@T�P ט ��T�T ��Q[R	 �BL�  �UCр D�*W[Q�_�_?ff�fe:lB ��P�ff@`�?33D  $a�U 3o>g�_�_po�l�P�e�9<�bbY���?٪``$o�oUAm��gD�`$�co�Quz9�P��Aa�P@a����C�Z`Ep�o]A63ffpu`aD/�U�h�͔r��~�a�R@ieAq�`�q��@9q�|�d&`%���c�333D�\P8���?�`?L�pAp[QB�b�k�}� ��z>�� >�ffԁL���T�f��fo � �Nw@�*�8�f���r� ,���П��ȟ��'�� ��F�`�J�X�����S�C�Vء��	�V3.00�Sl7r2c�T*��T�Q�� E����E�A E���E��3E��iNE�!hE��فEۑ�E��I�E��E����E�rF��F�F�M(F�5F�BFaOF��\F"f,�z�  E�@ E��� E�� E��  E����� �E����� E�ꆰԎ�ᆰ� �F   F� �F$ Fj` �F�@ F�P �F�` 9�IR/9�o���L�Q_ ��V���LQ�8TESTP�ARS�XUP9SH�Rk�ABLE 1%�J[4�SV�+�Q �0�V�V�VȨWQV�	V�
V��Vȥ�QV�V�8V�뱅�RDI��TQ�϶���������f�On߀ۊߜ߮�������Sl�RS 0ړ�� �����������#�5� G�Y�k�}��������� ����/]k�o��*	� %�7�I�����+�=��O؆�NUM  ��ETQ�P�P �밆�_CF�G ����Q@�<PIMEBF_T�Tq��RS~�;VE�R�<Q;R {1�J[
 8��RP� �@5  ������/ /&/8/J/\/n/�/�/ �/�/�/�/#?�/?Y?@4?F?\?j?|?{_��h@R
<PMI_�CHANG R >�3DBGLVQ`I�R;Q�0ETHE�RAD ?�E
;@�S �?�?TO6V��0ROUTe!�JZ!�D�OwLSN�MASK0HRSAA255.�E��O�O�8TOOLOFS_�DIq��5IOR�QCTRL �s[���n]8]_�_�_ �_�_�_�_�_o"o4o�Fo�
�_Tofo�og�PE_DETAIH�3ZPON_SVO�FF)_�cP_MOON �"P2�i�STRTCHK ��J^mO�bVT?COMPAT�h;C��d�`FPROG �%JZ%CAL�_TCP=�n%QP�LAYr��j_IN�ST_M�@ �|��g�tUSe]orL�CK��{QUIC�KME�0)�orSC�REF�3Jtps��or�a�f���2w�_{���ZyIS�R_GRP 1ξJY ؛  6�����;�)�_�M��8����Y�� �����͕�����/� �S�A�w�e������� ѯ�������=�+��M�s�	1234�5678����f�X�`�1�Ћ
 �}�ipnl/۰g?en.htm������0�B�X�P�anel setupF�}<�ϘϪ������� u�k�� *�<�N�`�r��ϖ�� ����������ߝ� J�\�n�����I� ?������"�4�F��� j�������������� _�q�0BTfx ������ �>�bt����3�~UALR�M�pG ?J[
  �*/!/R/ E/v/i/�/�/�/�/�/��/�/??<?�SEoV  �n6��ECFG ���m�6��A�1   ;Bȩt
 =?�s 3E�?�?�?OO+O=O�OOaOsO�O�Gz1ʂ҆�k SΟ�OH7I2sv?}{�`(%0?"_ p_I_4_m_X_�_|_ �_�_�_�_�_o�_3o��L� �M�OAoI�_E�HIST 1}��i  (p� ��,/SO�FTPART/G�ENLINK?c�urrent=e�ditpage,�t,1}o�o'{�(�o�emenu�b955�`�ou��(:L148,2 _XYd��` ����}_r_Z�������2�'C�M~69n�o� ��$�6�ŏN׏,68n��`4�@������3�M��}3�q���	��-���J���71n�MVn�������í�)a�a)o��� %�7�I�ȓޯs����� ����Ϳ\����'� 9�K�ڿoρϓϥϷ� ��X�j����#�5�G� Y���}ߏߡ߳����� f�����1�C�U��� �ߋ���������Я 	��-�?�Q�c�u�x� �������������� );M_q �� �����%7 I[m��� ����!/3/E/W/ i/{/�//�/�/�/�/ �/?��/?A?S?e?w? �?�?�/�?�?�?�?O O�?=OOOaOsO�O�O &O�O�O�O�O__'_ �OK_]_o_�_�_�_4_ �_�_�_�_o#o�_Go Yoko}o�o�o�oBo�o �o�o1?�og y�����o�� 	��-�?��c�u��� ������L�^���� )�;�M�܏q������� ��˟Z����%�7� I�؟��������ǯ ٯh����!�3�E�W��Bz�$UI_PA�NEDATA 1��������  	�}�  frh/cg�tp/wided?ev.stmc����ҿ����)  ri��.�Ip��F�X�j� |ώϠ�ϲ��Ͻ��� ���0��T�;�xߊ� q߮ߕ��������Bv���  �  - ��� @�E�W�i�{����� ��6�������/�A� ��e�w�^��������� ������+O6 s�l�� ��� ������1C �g������ �L	///?/&/c/ u/\/�/�/�/�/�/�/ �/?�/;?M?���? �?�?�?�?�?0?Ot %O7OIO[OmOO�O�? �O�O�O�O�O_�O3_ _W_i_P_�_t_�_�_ �_�_Z?l?o/oAoSo eowo�_�o�o O�o�o �o+�oO6s �l������ �'�9� �]�D����_ o�oɏۏ����#� v�G��ok�}������� ş,�������C� U�<�y�`�������ӯ ����ޯ�-�����c� u�����������T� ��)�;�M�_�q�ؿ ��|ϹϠ�������� ��7�I�0�m�Tߑߣ� ����:�L����!�3� E�W��{�� ϱ��� �������r�/��S� e�L���p��������� �� =$a����}�r�����)�*��V hz����� ���.//R/9/v/ �/o/�/�/�/�/�/?��������$UI_�PANELINK� 1����  �  ���}1234567890_?q?�? �?�?�?�4��]?�?�? OO1OCO�?gOyO�O �O�O�OYIY0:�M���[0  SOF�TPART/GE�NA1?CONFI�G=SINGLE�&PRIM=mainedit �O�I_[_m_YJ_$_M=�wintpe,1 @_�_�_�_�]�_$o6o HoZolooo�o�o�o �o�o�o�o
2DV hz����� ���.�@�R�d�v� �� �����Џ���~�M 0,  9P E=Por?S�5�co:�{�^������� ͟ߟ��'�9�� ]�o�R����O�O���� �Z1�/�%�7�I�[� m�`C�������Ϳ߿ 񿀿�'�9�K�]�o� �L���э͙�S���� �������#ߒS;�M� _�q߃ߕߧ�6����� ����%��I�[�m� ���2��������� �!�3���W�i�{��� ����@������� /��Sew��� �.���|�# G*k}`��� ���/�1/C/֤ �͡�ۯ}����/�/�/ �/�/?�2?D?V?h? z?�??�?�?�?�?�? 
OO�ϝϯ�dOvO�O �O�O�OE�O�O__ *_<_N_�Or_�_�_�_ �_�_[_�_oo&o8o Jo�_no�o�o�o�o�o �oio�o"4FX �o|�����e ���0�B�T�f�� ��/���������ُ ���>�P�3�t���i� ����Ο��O/�s/(� �/L�^�p��������� �?ܯ� ��$�6�ů Z�l�~�������#O5O GO�� �2�D�V�h� ��Ϟϰ�������u� 
��.�@�R�d�v�� �߬߾������߃�� *�<�N�`�r���� �����������&�8� J�\�n���������� ������m�"4ßX jM�q���� ��BT7x ������A��/ /,/>/P/C�t/�/�/ �/�/�/�/o/??(? :?L?^?Ϳ߿�?�? �?�?�? OO�?6OHO ZOlO~O�OO�O�O�O �O�O_�O2_D_V_h_ z_�_�_-_�_�_�_�_ 
oo�_@oRodovo�o �o)o�o�o�o�o *�oN`r��� ��m��&�8� �\�n�Q���u���ȏ ������"���?�?��{��$UI_P�OSTYPE  ��5� �	k�{��_QU�ICKMEN  ���j�����RESTORE 1ו5�  ���/
�2�D�h�m c�������¯ԯw��� 
��.�@��d�v��� ����W���˿ݿO�� *�<�N�`�τϖϨ� �����ρ���&�8� J���W�i�{��϶��� �����ߡ�"�4�F�X� j���������� �����y�+�T�f�x� ����?��������� ��,>Pbt�� ����( �L^p���I���� //��SC�REܐ?��u1sc-�uU2M$3M$4M$5M$�6M$7M$8M!��UGSER/ 4/F"T. �O#ksW#�$4�$5*�$6�$7�$8�!���NDO_CFG �؜�  ,� ���PDATE ��)�Non�e V��SEUFRAME  
���&,1RTOL_�ABRT7?��N3E�NBX?I8GRP �1�!��Cz  A��3�1��?�?�?�?�?FO"OG:�ېUx81g;MSKG  {5�Ag;N41%a��B%��O���VISCAND_wMAXyEI�c8��@FAIL_IM)Gy@f���#�8�@�IMREGNUMryG
�KRSIZyC�,���$,SO�NTMOUW0{D��%�VU�#�c�� �P�2F�R:\�O � �MC:\XS\wLOG�VB@4 !�O�_�Q�_o
��z MCV��_�SUD10fE�X9k
�f�wV�2�ꜙ�p(��=��͓o��j�o�o�o �o�o�o�o 2D�Vhz��KPO6�4_?S�0��n6�uQ0LI Q�z�xr�qV� �|f@�w��� =	�xSZ�V�~����wWA�I��DSTAT ܛ;�@�_ď֏��$����EP12D�WP  ��P G/����q�AP-���B_JMPERRw 1ݜ�
  � �2345678901�������ʟ�� ϟ��$��H�;�l��_�q����LT@MLO�W���P�@�P_TI�_X�('�@MPH?ASE  53���CSHIFT�UB1~k
 < ���Ob��A�g���w� ��ֿ��������� T�+�=ϊ�a�s��ϗ� ���������>��'��t�K�!��#ޛ:	�VSFT1�sV:�@M�� �5��4� �0��UA�  �B8���Ќ�0p������Ҫ��e@��ME*�{D�'���q��W&%�!�M�$�~k���9@�$~�TDINENDcXdHz�AOx@[O��aZ��S�︕��yE����G ����2�������<���RELE�y?�w�^_pVz�_ACT�IV���H��0A ���K��B#&��R�D�p��
1YBOX� ��-�����2�D�1�90.0.� 83v��254��2�p�&���robo�t�ԟ   �pN g�pc� �{�v�xx���$%ZABC�3�=,{�낆;- !/^/E/W/i/{/�/�/ �/�/�/?�/6??/?$l?!ZAT����