��   �S�A��*SYST�EM*��V7.7�077 2/6�/2013 A�   ����SBR_T  � | 	$SVM�TR_ID $�ROBOT9�$GRP_NUM<AXISQ6K �6NFF3 _PoARAMF	$��  ,$M~D SPD_LIT�  �$$CLA�SS  ������� � � VIRTUAL��' � 1 ��  �8���LR� Mate 20�0iC���BiSR1/60�00A��	H1 DSP1-� ���	P02.0�1,  	����PaR$� �� 8����M������
=����r��r����9"� �� ��� � ��� ?2� Er���  u�� �kk����� �Q��! 2�{(���=���4 �= ��c	1�����&�  5 ����� ��������� w���������2&�� �9�%�� 2 (�U_!N :?q�� T�/�/��/�/���/ ?�?%?7?I?��2�$����>�` ��( �H� 2�%�i0-��� �_ �C�>"�?�?�%72AzK�]o�8E"{;A��8r��퐵VT� $^����-��� � 1�4����?:�= �� � [l�q:��+
=� �� �r$ͥ?5$_ j?'5��M/_/q/�� �/T_f_x_�_�/�_��3�_�_�_o���@}�B> ��@wU�FBX'`X �oVo�4� "�?�10S.5�<=3AJ O�O n ��_c�K{n<D� �~��b
	QG�8CffH2e�� ~&$��?u3l���v�� �� � `���r�[�M� �����$�x]o5$� �?'���_  c/9	`R%Q��vx"���� �"�4�F��_j��_�� ����ď֏�������qo�e4/�5�m4A�a�oI@�a �b�d�R��ab1�k����m0��	z�{���t� 9 �7~��E���� 	��/���$�'�5#� d����5�|�����z¯ ԯ���S��?@�R��d�v�����������D)��e �11�h�5A2F����j��m�pq���h��.�.R�z3	y w�ݑ.g� ��������� � 3��� f�����5$��������!;��q��x"���(�r߄ߖߨߺ�� ��9���&�8�J�\�n�����B���76!��?9�K� ��`9H`.Y�qσ����9��ᶧϹς���  �q !����e	$���� �[7g"�݆Ss7� I�[�m�6HZl�� ��ߴ����� 2[7p����=UqQQ[7%v	v�ap� ����	//-/?/ Q/c/u/�/�/�/�/�/�/�/?<�?9?K? ]?o?�?�?�?�?�?�? �?�3oaO��� qO�O�O�O�O�O�O�O __%_7_I_[_m__ �_�_�_�_#?�_�_o !o3oEoWoio{o�o�o �?-OO�oCOUO/ ASew���� �����+�=�O� a�s��_������͏ߏ ���'�9�K�]��o ��u��o۟��� �#�5�G�Y�k�}��� ����ůׯ����� 1���U�g�y������� ��ӿ���	�ϗ��� 3ϭ���џ�ϫϽ��� ������)�;�M�_� q߃ߕߧ߹������� K��%�7�I�[�m�� ������#�U�G�� k�}�E�W�i�{����� ����������/ ASew���߭ ���+=O as�����)� ;�//'/9/K/]/o/ �/�/�/�/�/�/�/�/ ?#?5?G?Y?�}?�? �?�?�?�?�?�?OO 1OCO��[O��� �O�O�O�O	__-_?_ Q_c_u_�_�_�_�_�_ �_�_oos?;oMo_o qo�o�o�o�o�o�o�o KO}OoO8�O�Om �������� !�3�E�W�i�{����� ��ÏoՏ����/� A�S�e�w�������	 ҟş?Qc+�=�O� a�s���������ͯ߯ ���'�9�K�]�o� ��ݏ����ɿۿ��� �#�5�G�Y�k��ٟ �����!������� 1�C�U�g�yߋߝ߯� ��������	��-�?� ��c�u������� ������sϥϗ�`� ���ϕ����������� %7I[m ������G�� !3EWi{�� ���1���g�y� ��S/e/w/�/�/�/�/ �/�/�/??+?=?O? a?s?�?�?�?�?�? �?OO'O9OKO]OoO �O�O//�O%/7/I/ _#_5_G_Y_k_}_�_ �_�_�_�_�_�_oo 1oCoUogo�?�o�o�o �o�o�o�o	-? �O�O�O��O�O�� ����)�;�M�_� q���������ˏݏ� ��oo%�I�[�m�� ������ǟٟ���Y "�����{����� ��ïկ�����/� A�S�e�w��������� ѿ-�����+�=�O� a�sυϗϩϻ�7�)� ��M�_�q�9�K�]�o� �ߓߥ߷��������� �#�5�G�Y�k�}�� 뿳����������� 1�C�U�g������ϰ� ������	-? Qcu����� ��);��M q������� //%/��J/=/���� ���/�/�/�/�/�/? !?3?E?W?i?{?�?�? �?�?�?�?�?UO/O AOSOeOwO�O�O�O�O �O�O_/Q/�Ou/�/�/ a_s_�_�_�_�_�_�_ �_oo'o9oKo]ooo �o�o�o�oO�o�o�o #5GYk}� �O__�3_E_�� 1�C�U�g�y������� ��ӏ���	��-�?� Q�c��ou�������ϟ ����)�;�M�� r�e����˯ݯ� ��%�7�I�[�m�� ������ǿٿ���� !�}�E�W�i�{ύϟ� ����������߇�y� #ߝ������ߛ߭߿� ��������+�=�O� a�s��������� ;���'�9�K�]�o� ���������E�7�  [�m�5GYk}� ������ 1CUgy��� ����	//-/?/ Q/c/u/���/�/ +�/??)?;?M?_? q?�?�?�?�?�?�?�? OO%O7OIO�mOO �O�O�O�O�O�O�O_ !_3_�/�/K_�/�/�/ �_�_�_�_�_oo/o AoSoeowo�o�o�o�o �o�o�ocO+=O as������ ;_m___(��_�_]�o� ��������ɏۏ��� �#�5�G�Y�k�}��� ����ş����� 1�C�U�g�y������ ¯��/�A�S��-�?� Q�c�u���������Ͽ ����)�;�M�_� q�͟�ϧϹ������� ��%�7�I�[�ׯɯ s������������ !�3�E�W�i�{��� ������������/� ��S�e�w��������� ������cߕ߇�P �߽߅����� �'9K]o ������7�� /#/5/G/Y/k/}/�/ �/�/�/!�/�/Wi {C?U?g?y?�?�?�? �?�?�?�?	OO-O?O QOcOuO�O�O��O�O �O�O__)_;_M___ q_�_�/�/�_?'?9? oo%o7oIo[omoo �o�o�o�o�o�o�o !3EW�O{�� �������/� �_�_�_x��_�_���� я�����+�=�O� a�s���������͟ߟ ��_�9�K�]�o� ��������ɯۯ�I� �������k�}��� ����ſ׿����� 1�C�U�g�yϋϝϯ� �������	��-�?� Q�c�u߇ߙ߫�'�� ��=�O�a�)�;�M�_� q����������� ��%�7�I�[�m�� �ϣ����������� !3EW�����ߠ ������/ ASew���� ���//+/��=/ a/s/�/�/�/�/�/�/ �/??q:?-?�� ��?�?�?�?�?�?�? O#O5OGOYOkO}O�O �O�O�O�O�OE/__ 1_C_U_g_y_�_�_�_ �_�_O?A?�_e?w?�? Qocouo�o�o�o�o�o �o�o);M_ q���_��� ��%�7�I�[�m�� �_o�_ȏ#o5o��� !�3�E�W�i�{����� ��ß՟�����/� A�S��e��������� ѯ�����+�=��� b�U�Ϗ�󏻿Ϳ߿ ���'�9�K�]�o� �ϓϥϷ��������� �m�5�G�Y�k�}ߏ� �߳���������w�i� ����y���� ��������	��-�?� Q�c�u����������� +���);M_ q����5�'�� K�]�%7I[m �������/ !/3/E/W/i/{/���/ �/�/�/�/�/??/? A?S?e?��?}?�	 �?�?OO+O=OOO aOsO�O�O�O�O�O�O �O__'_9_�/]_o_ �_�_�_�_�_�_�_�_ o#o�?�?;o�?�?�? �o�o�o�o�o�o 1CUgy��� ����S_�-�?� Q�c�u���������Ϗ +o]oOo�so�oM�_� q���������˟ݟ� ��%�7�I�[�m�� �������ٯ���� !�3�E�W�i�{���� �����1�C���/� A�S�e�wωϛϭϿ� ��������+�=�O� a߽��ߗߩ߻����� ����'�9�K�ǿ�� c�ݿ���������� �#�5�G�Y�k�}��� ������������ {�CUgy��� ����S��w�@ ���u����� ��//)/;/M/_/ q/�/�/�/�/�/'�/ ??%?7?I?[?m?? �?�?�?�?�?GY k3OEOWOiO{O�O�O �O�O�O�O�O__/_ A_S_e_w_�_�/�_�_ �_�_�_oo+o=oOo aoso�?�?�oOO)O �o'9K]o �������� �#�5�G��_k�}��� ����ŏ׏����� {k