��   �A��*SYST�EM*��V7.7�0107 10�/3/2018 �A ���$$�CLASS  O���(��D���D VIRTUA�L%7MNUFR�AME AF�D� �� 	 88�?���}��y�� ����1= gQs�������	/�/?/��WN_UM  ��>lx�  WTOOLa�4 
wN%M/ 7 Bp�#C>3/U/ �/1/	?3????i?S>�$����D}�?:�1>�y]�1�1>Ӌ��&  G __?�?�? ]?�?OO%OOO9O[O��OoO�O�Og,�!{&
���&* 