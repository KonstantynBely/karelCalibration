��   3L�A��*SYST�EM*��V7.7�0107 10�/3/2018 A   ����UI_CON�FIG_T  �d )$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$DU�MMY37CME�M_LIMIR$DBGLVL��POPUP_MA�SK�zA  u�8�ODE�
]9CFOCA �[40CPS)C��g 
HAN� ~� TIMEOU��PIPESIZE{ � MWIN�PANEMAP� � � NU_F�AVB ?� 
$wHLP> _DIQ�?� mELEM�V}UR� h� S|o�$HMI��RO'XW AD�ONLY� �T�OUCH�PRO�OMMO?$��ALAR< �F�ILVEW�E�NB=!%bC �-"USER6)FC[TN6)WI�� I* _ED�h"R!�_TITL� ~-"COORDF8"}&USTOM0� t $} R?T_SPID��$�C�$*PAG� ?�ZDEVICE��)SCREqEF����'N�@$FwLAG�@  &�USRVI 1 O < \� �;2�<1PRI��m� A� [0TRI�P�"m�$$CL�ASS  �S��|1��R��Rq0VIRT_1z?�0'�2 )�U�)�_�pR	� �,��$;����2�0�3�3��1�� , ��  �?��
 ���1<ONO`OrO�O�O�O 8O�O�O�O __'_�OK_]_o_�_ �_�_4_�_�_�_�_o #o5o�_Yoko}o�o�o �oBo�o�o�o1 �oUgy���� P��	��-�?�� c�u���������L�Ꮐ���)�;�M� �TPTX��p݈p���  sX����$/soft�part/gen�link?hel�p=/md/tpmenu.dgO� �����؏C�U�g� y�����,���ӯ��� 	����,�Q�c�u��� ����:�Ͽ���Ϭ)���9���F�6�3S�($ÿ���� nϧϒ������1�1@���3a�Y��?����9�3�" 1�5�2� \�6 �REC VED���i�{�whol�emod.htm���singl���doub��t�rip��brows��+�|��0� B��f�x�������f�P�ߜ�dev.Es��l$���<�1'�	tS���<��� ��� ���������� 2[� �0s�� ����� 0pEW&{�� �]�VP���/ /,/>/P/b/t/�/�/ �/�/�/�/�/??�� .?(?V?h?z?�?�?�? �?�?�?�?
OO.O@O ROdOvO�O�Oh�O�O �O__/_A_S_e_w_ r�_�_|_�_�_�_� ��O=o8oJo\o�o�o �o�o�o�o�o�o "4]Xj8?�� �������0� B�T�f�x��������� ҏ����O1�C�U�g� y���������ӟ�_�� 	�؟�?�Q�oo � ���������ܯ� � )�$�6�H�q�l�~��� ����ƿ���� � 2�D�V�h�zόϞϰ� ��������
��.�@� R� ��ߟ߱������� ����/�*�S�e�4� F���d�v�\����� ��=�8�J�\����� ������������ "�B<j|�� �����0 BTfx���|� ��//1/C/U/g/ y/�/��/�/�/�/�/�	?:�$UI_U�SERVIEW �1��R 
���J?\?�m{?�?�?�?�? �?�?O"O4OFOXO�? |O�O�O�O�Oo?�O�O �OgO0_B_T_f_x__ �_�_�_�_�_�_�_o ,o>oPobo_oo�o�o o�o�o�o�o: L^p�%��� ���o����C� l�~�������W�؏� ��� �ÏD�V�h�z� ��7�������/���
� �.�@��d�v����� ����a������*� ՟7�I�[�ͯ������ ̿޿����&�8�J� �nπϒϤ϶�a�k� ����Y��4�F�X�j� |�ߠ߲������ߋ� ��0�B�T���a�s� ��������������� ,�>�P�b�t���)��� ������������# ��^p���I� �� �6HZ l~)3��!� �/ /2/D/�h/z/ �/�/�/S/�/�/�/
? ?�(