��  ë�A��*SYST�EM*��V7.7�077 2/6�/2013 A�Q  �����ABSPOS_G�RP_T   � $PARA�M  �  �ALRM_�RECOV1   $ALMO�ENB��]ON�iI M_IF1� D $ENA�BLE k LA�ST_^  d�U�K}MAX�� $LDEBU�G@  
GPCOUPLED1� $[PP_P�ROCES0 Ľ �1����UR�EQ1 � �$SOFT; T_�ID�TOTAL7_EQ� $,�NO/PS_SP�I_INDE���$DX�SCRE�EN_NAME ��SIGN�j��&PK_�FI� 	$T�HKY�PANE�7  	$DU_MMY12� ��3�4�GRG_�STR1 � �$TIT�$I��1&�$��$�$5&6&7*&8&9'0''@�%!'�%5'1?'U1I'1S'1]'2h"�GSBN_CFG�1  8 $�CNV_JNT_�* �DATA_C�MNT�!$FL�AGSL*CHE�CK��AT_C�ELLSETUP�  P� HO�ME_IO� }%:3MACROF2�REPRO8�DR�UNCD�i2SM�p5H UTOBAC�KU0 � ��	DEVIC#T�Ih�$DFD��ST�0B 3$�INTERVAL��DISP_UNsIT��0_DO�6�ERR�9FR_F�a�INGRE5S�!Y0Q_�3t4C_WA�4�12HG�X_D�#	 d� $CARD_�EXIST�$�FSSB_TYP�i� CHKBD_[SE�5AGN G�� $SLOT�_NUMZ�APR�EV��G �1_�EDIT1
 �� h1G=H0S<?@f%$EPYO$OPc �0LETE_OKzB{US�P_CRyA�$�4�FAZ0LACIwY1KR�@k ~�1COMMENy@$DGV]QP�� ���AL*OU~�B , $�1HV1AB0~ OLz�UR"2CAM_;�1 x�f$�ATTR��@0A�NN�@�IMG_�HEIGHyAcWoIDTH�VTC�YU�0F_ASP�ECyA$M@E�XP;$� Mf��CFcD X '$GR� � S!1U`=BfPNFLIC`~d
UIREs3��A�OMqWITCH�}cX`N.0S_d�SG�0 � 
$WARNM'@f��@�� LI? �aNST�� CORN��1F�LTR�eTRAT�@0T�`  $ACC�1"p '|��'rORIkP�C�kR�Tq0_SF� �!C�HGI1 �[ Tz`u3IPpT�YVD�@*2 �P`�`� 1zB*HD�SQJ* ��q2�v3�vU4�v5�v6�v7�vU8�v9��vqO�$ <� so�o�h�|s1�PO_MOR.� t 0E�v�NG�8`TBA� 5c���A������]@����ϋP��0Ѕ*��h�`�
P�@�2� �,p�J�,p_Rrrqo@+�J�/r/�J�JVq@�C�j��m�g��ustP_�}0OF� 2  @�� RO_���WaIyT8C��NOM_�0��1ەq3W ��cDC �;����hP����mEXpG�0� xF�p%r
$TFx�lJF�D3ԐTO�3�&@U=0�� ��H�24�T1��E�� �e��f��f|��0CPDBG;a�� k@$�PPU8�3�f):��&A�AX 1�dUN�$;AI�3BUFuF����! |�`��`[PI��Pr�EMq�M~�䠁�Fr�SIMQS��G�h�QE�����MC{�k �$}1JB�`S�}1DEC�������۵z� ě0CH�NS_EMP�r#$Gg�=Ǎ@_��q3�
p1_FP󔞡TCh�@`�b��q0�c}�y�G�� V�AԂ�!!���JR!0ԂSEGGFRA.pv 7aR��T_LIN�C��PCVF������Y ���Q��)B����( '���f�e �S���Q��.0�p�B�8�A����SIZC����z�T��g������QRSINF3��p�� ��?�������؉����Lot��G�*�CRC�eFCCC�`+���T� h��mh�SbA��h�*��f��:�D�d�c��C��PTA����w@��L����EV���jF��_��F��N&�G�� �X������1i��! ��,��h#RGNP��0qF���R�}�D���2}�LEW N��Hc6���C�K�|A�dCx :�@L��ou2���A6N`�Co�$LGp��B@�1aP��s@�dWaA?@����~0R���dM�E%`��d�_RAs3dAZC���z��OkqFC�RH`X`F�`��}��,�ADI ;� 6b� ���` �p�`5cn�S�@1�L7a�AMP���PY8C�U�MwpU��iQU� $�P��C�C�G1������DBP�XWO����p�$SK��2��DB]T TRL�1 ���Q0Ti� �P�DJ��4LAY_CAL`�1R !'PL	3&@�0ED�Q5'�Q5'"̡���1!�W�;PR� 
�1� 0�1" �PA�$�q$�� ��L�)#�/�#mp�0$��/�$C�!%�/���2PEqr�&�/�#�d REp�"'H� �O)@"$LF3#$�#xB� W;4���FO[ _D0m�RO(@���u��j��~�3RIGGER�6�PA%S���ETUsRN�2RcMR_���TU�`?�u0EW5M����GN�P���zBLA��E��$�$P#�CP� ��&�@�Qk�C5D�mpD��A#�p4\1i�FGO�_AWAY�2MO���fQg�CS_n(<�QIS  ����c�C���A����B�t�Cn��A"r�FW���DNTV@��BVkQ�����S˳W��sU�J&�U�� ��S�AFE�ZV_SV>6bEXCLUl������ONLA��SY���Q�tOTBa��H�I_V/M�PPL�Y_�a��VRFY�_#�q�Bd�_ #)0���_+�Ipg `"�@SG3� *�b݀�0 AM�@��a*����0��Vi|.b%fANNUN� ,rLdIDp�U�2~S@�`mijarj�f�(�堫@I�"+��c$FOb�׀OT@�w1 $DUM�MY���d[!�d١��& �E, ` 8�HExs��b�S|B$�SUFFI��@ ��@�a5��g6�a��DMSW�E- 88�KEYI����TMZ1^ӌqL�1�vIN������. D��HOST? !�r���t�[ �t٠�tYp�pEMp>���$��SBL��;UL��/ �|�3����T50�!0 ϴ $9��ESAMP�ԕF���������I�0��$SUBe�Q�� �C�:��G�SAV��r����G�C� ˇ�PnfP$�80E��YN_Bn�1 0�`DIadb�@O���}$]��R_I�� �E�NC2_ST � 2
ԇ J���L�q~S�`;����!3�M�I��1:�p�4  AL�3�M��0�0K�4x'a��AVER�q8��}�M�DSP�v��PC�U���\�ެ�VALUŗHE4� ��M�IP@����OPP7  �THS ���6�S�F�	F􁳠dL�0�T���SC�Q�d:�ET�o�5zrFULL_DUY�da�0��O�w�h�OT���0�NOAUTO�!6��p$�\���cTl�
�C` �C����`!�L�� _7H *�L���n�b���$�0P�˴ ��ֲ��[!���a��Yq���dq��7��8��9R��0����1��1��U1��1Ⱥ1պ1�U1�1��2
�2�����2��2��2Ⱥ2�պ2�2�2��3J
�3��3����3��U3Ⱥ3պ3�3��3��4
²q��SE�"8 <��~��`��;I�����/��QFqE�0�0� 9 ,���Q? z@^ ?Q�А��ER@�#�`!�A��� :�`�$TP�$VA�RI�<��UP2f�P; �pq�TD�� �S|�1`3���qr�wBAC�< T�pr��)��bP�P o�IFI)�P ���U����P��*��F�0��� =t �;'�Ԡ��P'�ST (&�� HR&�r0E��*��	%�C��	��� _Cr�N�r��B��p�h�FORCEUP%b^n�FLUS�`H�N �E�h�RD_C�MK@E(����IN�_��&vPg�REMM�F~Q��M �� �3
K	N0�EcFF��N@IN�A��OVMl	OVA�l	TROV���DyT��mDTMX� ��m{@�
��? �*X[ ��CL��_:p�']@$�-	_
�;_QT��X
��@AQ	D� ��}��}!�V1� RQ��LI�MIT_�a椀�M���CLmd}�RIqV	�a��EAR��IO*PCC�����B�Bg�CM@��R{ �GCLF��G!DYM(/�aR#5TWDG��| s%� �SS& �s> �P�a�!r1��wP_(�!�(�!1��E�3�!�3�+5�&�GRA����?w��kPW晅ONT��EBU�G)S&2*�P{@a�_/E @�P�Q�`_�TERMB5AK5N�QORIG0BK5�`�SM_�Pr�G0�Cd9TA�9Dd6� �UPB�E�3 -zAa�@.PY3>.@A$SEG�:f �ELEUUSE�@NFI,��2�1ޠ<p4�4B$UF6P��$�FQ4@��wAG0TQ�&�HSN;ST PATm�p�iBPTHJ�AߠE �p��2�P؀	E)�؁���1R�@�InaSH�FT_��1oA�H_SGHOR ܣ�6 �0�$�7�@Dq�'�OV�R#�na�@I�@�Uz�b �QAYLO=�z��I'"�oAj�!�j�ERV��:Qh��J ��OG @�B0����U>����R!P"�ASY1M.�"��1WJG�т�ES�A�YvR�U��T @���E)�ᥳEP�!�WP!�WOR @M|B��GRSMT��F�GR��3laP�A.@��`�q�uG ׸ ����TO�C�1�`P�@ �$OP��ဝpՓá �e�O��RE�`�RC�AO�pтpBe�`RmE u�h�A���e$PWR�IM�ekRR_�c4��qB� H2H���p_�ADDR��H_LENGqByqnq�q�uR��S�I H��S���q0Ӧu>Ӵu����u��SE�'�LrS<��J $N�`���_OFF��rP�RM� ^�aTTP_�H�wK (^pOBJ?"lip��$��LE`C�!�ȠL � \�׬�AB_~TS�bs�S{`��*�LVN�sKR��eHIT��[BG��LO�qt��fN�͂���`���`SS{ ��HW��A��M�p`INCP}U�"VISIO� ����+��t,��t,���� �IOLN��N�̠�C��$S�LQb��PUT_&�$�`{�P ��V���F_AS�"O��$L��I����A"��U�0�@Af��`q�<PHY���ÓZ�析UO��#P ` ������ڔ� �2�pP���`(�L��Y�,B�Z�UJ�Q�z�;NEWJOG-G���DISx�SV�K�-�f�#R 
�WAV��ǢCTR�CǢFgLAG�"[�LG�d�S ���Y�3LG_SIZo����������FD)�I �4�E�*��D0�� �c$���𖶦���K��D0��� SCH_ ��߅p�2��N��F�T���E�"~���D����U
�
�{`L�n	�DAU/�EA��-��dE�;�GH�b }��OGBOO��Uh Aɒ��I�T��y�[0ŖREC���SCR��ʑDeIēS.@��RGO� ��˒����d�´���	SU���W�Ĳ�Ľ��JGM$�MNCH|,�FNKEY%��KM�PRGK�UF�Y�PY�FWDY�H]L��STPY�VYذ@Y؀�Y�RS��H1`uۺ�CT���R��� �$�U	�m���
R��ݠғ`�G=��@P�Od�ڻŦ�M�F�OCUd�RGEX.��TUIK�I{�����	������I�M��@A�S�`���@������ANA���2�oVAILl�CL!~�UDCS_HI+4�`�s_�Oe�
!h�SȚ��|�S����IGAN4��F�J��T�bL�8�BUj � V 5!PT�$*���rv�Ϥl1��AVrW !Pi�'���0�1?2?3?_�>� X � i�=a0�5���Ņ�ID� tb	P5R�bOh ��\A�+ST	�RF�Y� �@~�  W$E�C�y�����!���!Y L�؟0� �@���`qFtǀ�Fw�Ҭ�_ Z �i`����b���>0C���[ �p CLD�P	��UTRQLI�{��T����FLG �� 1�O�D������LD���ORG������hW>(�spiT�r� 4\ �#0P��վ�Sy`T��70#0' �$�!�#RCLMC�$B/T/�)�Q��!=1I�p_d] �d�RQ73$DgSTB�p�   6l��-8AX�R /8�I<EXCES�bR 5Mp�1^��2��T2��0_�p"6_A:&��;G?Y8�0K�d` \�G�ROU��t$MB� �LI9�CREQGUIRDB�aLO#KODEBUr� 1LYM��agbʑ`@�C�"MND��`c`ab���̨�CDC���IN'��C��Z`����H��N��a#�� �EPST�� cn\rLOC�RITp��P�Ap�1 1�ODAQ��d X&�ON�cF�R� fV�	X��b�U���u�u�FX0IGG>�� e �y X��a��X�XR�Q%��Y	��X	��V�0�ғDATA$`E��a��a�N��f �t $MDEaI�:�)Sf��^d�![gH�5P�@]ez��a_cAN�SW�a^d�a��^eD��)ARz�� Xpg -�0CU4�V�`��=URR2{�h D�2�`A��A�! d�$CALI&0��GtS�w2K�RINb�:t<�NTEg�(�i�bCu��=RBqg�_N�qjPukr���$ht��2kuyDIV�&D�Hi0jp+�l $�Vp�C�$M��$Z0R<!T 0R����b�emH �$�BELT˪ZACCEL���;�"��IRCO�݁m��T<���$PSi0�Lt�ڰW��Cp8�x�T�9�PATH����.���3]��Pl1_@<�r��Ł�"S Cr���_MG��$D�D�9���$FW��`7`���.���D}E�PPABNe�ROTSPEEՂ@L� JN�@��(0��t�$USE_dp�P&�ܦSY>���p�! �QYN0A�����OFFua��M�OU߁NGJ�܀O9L~�ٔINC�d2Q���-2��� -2ENCSpa2U��+4R�IN�I��B�����"n�VE��s^�2�3_UPօp�LOWL��[�` '���D>�2@Ep]'�r�2C[pW�MOS����4MO��0�'PE�RCH  ��OV ����蓼������$ �8S+�� 2@������!V�0^�O�L�P��7O�U�UP"�����Ω�TRK��AYLOA�J��1�����͵³3P� �RTI�1	�� MO�O�-2@�28 �`4�wٳx��?�pDUM2���S_BCKLSH_C��P�ϐΦ�����bn�"�y�Ñ��!CLAL V��!��� N��CHK �SՐRTY����C�
*!r6a_�ä_UM��r��C���SCL��W�LMT_J1_�L< 0-օa:�E�4�U�G�D�J�P�J�S�PCd�ȑZ���3�P	C �3�H_A@��řC� cXT���C�N_rN���.�S��%�V���:����ѹ�9���C' �SH�r�*�*!9�9�� p��^���9���PAL���_P��_��"�Ŷ�!ճ����J1G����~�OG��,��TORQU��ON ��޹*�B٢-�*�L�_Wž�_�sj��s�j��sj�Ir�I��I�sFKP]�J�!��c!�VC�0'4�2���1��{0��82��JR�K��+� DBL�_SM���"M�@_sDL�q�"GRVq�`j�sj�sKH_��8I���
COS���LN- �����p �	�p�	�����F1Z� ٦KMY�D�TH�eTHE{T0��NK23�s؏�s� CB�CB�sC&1n2�����s���SB�s��GTS�1W�C.�2Q������$�'3$DU���8A!r��2�P&��1Qb8V$N	E�4�PI� ���"%�v$�p�A��%�'8���LPH�5�"h��"S��3�33@�"+3:2�pV�(QV�(�p�,V�*V;UV;V";V0;V>;VL9H�(�&�2�-n�TH;H;H";H0;UH>;HL9O�,O�(�O}I�.O�*O;O�;O";O0;O>;O2F�"�Y�T�'�SPBALANC�E_T@SLE�H_�SPHq�hR�|hR3PFULClX`�R{W�R3Uz1i
��UTO_����T13T2�Y�2N��� `��Tq���Ps d����T�O�p!�L�I�NSEG���REqVf��Q�DIF��fzy1j_g�r1k���OBUa��t$yMI�`���SLCHWA�R>��AB��u$MECH�Tˑ,�a��AX˱Py��f8�'�r�Pl 
�bI���:�ROB�CR�W�-u���*�M�SK_KP�tn P+ �P_��R��r_tn���18�c�a�_p�`�y�_p�aIN:a��MTCOM_C|���po  ݀�g`4�$NORE�S��r��`�rp �8U�GRJ��eSD�� ABג$XY�Z_DA�!F�r�D�EBU:a�q���pqu _P$��COD��G 1����`���$BUFIND�Xa�  !�MO�RRsr $�qU@&���u��ӑy�^���bGi�s � ?$SIMUL��8���>���F�OBJE|jP��ADJUSψ�AY_I��8�Dp���s�Ԑ_FIב=s�TZ��c�� ��`b�"�(�b`p0G��D��FRIW�d�T&g�RO%�A�Eb�=^�OPWO> Vp�t0>�SYSByU0[�$SOP���I�����U��b`PR�UN�rڕPArpDpٖ�b��1�_OUT�Α�a�t$�I�MAG��\pv PfDaIM��1�IN[ ��0�RGOVRDY�˒���P�/�a�� L_�PB�}����SRB�� ��Mkᦜ�EDb��` �N2�@M��~�SW��]��SLjPVpu x �$OVSLfS;DI��DEX���q �����o��Vb��N�A��'��,�'��D�M~]�ӣ_SE9TK�Vpv @U�^�L�ep�RI��j�
q�_�}�����Z�dà>*� w H\q�`���ATUS<�$�TRCx T�X�ѳBSTMڷıI��P��4}Ѱ���Vpx DB\pE���β�0Ehb�ϱ�����ϱEXE�հ����)�=��f�y�m�]p԰UP�L�9$�`6�XNN����x������ �PG�u7zWUBñ�e���ñ��JMPWAeI[�P���LO7���pFA`��$RCVFAIL_Cwq�p��R9��p�c��(��}�"�-�AR_PL��DBTB��,��pgBWD ��pUM*��"�IG�7��Qc�T#NLW�"�}�Ry�iӂ��E�����^���D�EFSP` {# L\p�`��_��Ճ��UNI����Ѐ��RD��Rb _LA`PFͱ�ѦpUq|-��#��q�O��XPc�NN�PKET�
��Pq�Uq} h�ARSIZE5p��=���u�S̀OR��F�ORMAT�Pg�C�Oנq�<bEM�dL����UX��,����LIb�Uq~  �$�pP_SWI��`��6^�/ G�b�A�L_ o���AR�rB���C�rD���$EL���C�_lі� � �c ���r��J30 ��r��TIA4Z�5:Z�6�rMOM��f��s���pB��A�Df��s����PU�NR����s����������Rt�� A$PI�&E�kqE�p -~-�-�WC �0$��&�9q�g|E��eSPEEDL@G�����Ծ���� )�9����)��	)���SAMWPx�0�1��MOVD�H$_@S`Y%nk%_��1�t�2�t����c�v��28�H�PxIN��� ������(�<+(+GAMM<Vu!>�$GETE�U��ٓD5�
�PLI�BRv���I�$H�Iu�_L�ݰpB�&E��(A�.� �&LW �-�&�,�)	6�&1��f��`j��� $�PDCK���ٓ_�����E����b7��a4��a9�� �$I��R�`D`�c�b~�Ե`LE�q`kq���81��0���ܑ`Vp�P/aUR_SCR��A�r���S_SAVE_DX��8Ex�NO5�C�� y�6�8@{$E�.{I�� G	{I�@�J�KP�q� �H� ���x"Mao ���s����d���6W2U�Cqy����M� �k�F��a�E��3�W<�@[�jQWg@5r�U�R�R��Sdc2jQM"��[CL�W���M)ATr� � �$PY����$W`�fNG�O�` �b�b�b#�H�@���a� ���c��X�	O���Z�e��ހRtG� p䠰p�3+�zO�O�O�O�O�a5�_�r� |�E�8@�� >vs�>v��8@_�kwVv�y�Eހu%X� tB��\�P�"tP���P�M&�QU5 �{ 8*�QCOU�1� �QTH#pHOL�<�QHYS��ES�e�qUE�p.BZ�O.��  q�P���%杲UNְ�Q r��OE��p� P2��3��AÔ�ROG(�����Q2(�O}�2�x�����INFO�q�� #�e����R�v��OI��� (�0SLEQ�с�рHi�C�{�D��L��`�� OK0r��!E�� NU!��AUT<TA�COPYqu�(?��`@ML�NI�M��X�Cᐛ� Y�RGWADJ�q�i�X�Q���$ഖ�`��W��P���0�������[EX8�YC0b�ђ�Obp�q���$�_NA9!��������`��� � 9Q���POR�A�\B�SRV0�)a�6Y�DI��T_��{��������������5*��6��7��8y����S8BL��m�MC_)F�p��PL9A8An�ȰR��9��Ѽ���$iB����d� ,ƨ0FL-`L�C@YN��[�M��C?��P�WRc��L��!�D�ELA��8Y5�A�D�a��QSK;IP� �Q�4�-OR`NT�Q ��P_4��ַ@lbYp �������� ��Ƞ��ՠ������z��9�1�J2R� nL�� 4*�EXs TQ%����(Q�����p�����p���RDCNf� �`��X9�R�p�����r��A$�RGEAR_� I9OT�2FLG��vi̥�M%PC��B�UM�_����J2TH2yN'�� 1������G8 T00 �$����MlѺ`I�8��qREFr1�q�� l�h��ENAB{�(cTPE�0�1� ���i�m���^QB#��@:��"������2�������������&�3�Қ7�I�[�m����&�4�қ������P�����&�5�Ҝ1�@C�U�g�y���&�6�������������&�7�Ҟ+=Oas�&�8�ҟ������&�SMSKJ�q�|��a��E?Aި�MOTEF�����a@��(Q�IIOQ5�Ic(P���POW�0L�� ��pZ����#p%�L���U�"$DSB_S�IGN�1)Q%���C�l�(P���S232���b�iDEVI�CEUS�,R'RP�ARIT��D!OP�BIT`QY�OWCONTR;�(Q�ѬO'RCU� MDSU_XTASKT3N�p�[0�$TATU`P#6V"�0L����p�_,PC9�$FREEFROMSp���%�GET�0�U�PD(�A�2V"P|� J��� !)$USA^���6<���ERIO�P@&bpRY�5:"_>@ �qP}1�!�6WRKI�[D���6��aFR�IENDmQ�P$�UFw���0TOO�LFMY�t$L�ENGTH_VT�l�FIR�`-C�RSyEN ;IUFINR:]��RGI�1ӐOAITI��4GXӱlCI�FG2�7G1�0�Ѐ3�B�GPR� A��O_~ +0!�1R�EЀ�E3�e�TCp���Q�AV �G8��"J���u1~! � �J�8�%��%m��5�|0G4�X _0*)�L|�T�3H6��8P���%r4E3GU�W�P�W�R�TD����T���а��Q�Tm�$V 2����1��R�91�8�02�;2/k3�;3�:iva�9=i��aa�^S�jR$V��SBV�EV'�V�B
K�����&c�p���F�"{�@�2q�PS�E��$.rRC���o$AŠFwPR��Gv]U�cS'�� 7�sA6I�� 0�@DqV`��p�d`���PE0�@��=�
B5S!/� ��aRg�����R�6�N AX�!$�A�0L(A���r/THIC�1Y���h�t1TFEI��q�u�IF_CH�3�qI0�G�a�pG1bxf�з�m���S@��_J�F��PR�ֱ�S���Ԁ�d �$�SР�Z�GROU��̃TOT�t̃D;SP�JOG���#&��_P��"O������j��&KEP(�I�R����@M�R@�A	P�Qn�E^�`�!�[��SYS6��"[�PGu�BRK�B �.��pIq�p��M���΂��`AD�!̃9�BS�OC׆�NӕDU�MMY14�p@S}V�PDE_OP�#�SFSPD_OVR=���C����OR�CNm0�F�.����OV��SFR��pU���Fn��!#�p�C��A�"LCH�����РOV�s0��Wb�@M��ĥ:�RO�#�ߑ�_�p�� @�@�u@VER�ps0O�FSu@CV? �2WD6���2�ߑj2Y����TR�!���E_�FDOY�MB_CiM�D�B�BL�b>�f��attV"Q�240�/p��N�Gg�z�AM�x�Z�0���¿_M�~��"7����8$C�A�7�D����HcBK81��IO�5q���QPPAʀ=�"�M�5�͵���DVC_DBxC~� � 3"�Т�!��1�����3����pН�*���U�3��CAB ��2VӆPѣIP��c��O��UX�SUB'CPU�r	�S�P  P���90^SQ׹c��."~��$HW_C�А���S��cA�A�pl_$UNIT��l��ATTRI"���	��CYCL��NEC�A��J�FLTR_2_FI_�G(��9&��1LP�?�>�_S�CT�CF_��F_��6��FS8!����CHA�1�wᇲ�"v�RSD�4"�����q�_T��PROX��>�� EMy_ܠr��8d��a d���a��DIb0!�RAOILAC��9RM��CLOÐ C��Q*q���3q���PR��S�Q�pU�Cr�� 	��FUNC��@rRIN'PѸ0��u��!3RA��B ����8F�Ğ�WAR~���#BLQ����A��������DA����	����LD)0��Q1�q2��*q1TI2rQ�ǁ�p$xPRIA�1�"AFB�PP!�|ߠ�<`�R���MsOI��A�DF_&@؅�51��LM��FAށ@HRDY�4ORG6 H���A�0 �MULSE&@"�Q��a �G�	���m��$d$�1$1 ���0��߮� xm�EG0�̃�`ARހ���09�2o��z�A�XE�ROB�Wd�A��_�œSY������S�WRI�@s1��STR��� ��(�E�� !	%1��AB( �/&�a�ӰOT0v^�	$ߠARY�s�f"���S@	�FI���*�$LINK(���!�a_%#��%{q�"XYZp82�*�q�#OFF��R�"�"�(j Bဂj�4С��n�3FI��%7�q���j����_J���%��#�QO�P_>$H+5�3�PT�B\1�2C��i�D�U�&62�TURN��2r�5t!}��p��|7FL�`���m�0��%+*7�	� 1��. K�M�&8�2�Q�2rQ�#�ORQ ��G��-(�+p��z��� 3q�E"��T�GOV�@-A��M*�y�4 �E:�E@�FW�J� �G���D��o�*� � �A7�P��y��E�A�G`ZU:ZU�CG�ER�
��	6�E���B�TAFQ��)4����r'�AXУa2.q �c�W�c�W�c�W�p�Z �0�Z�0�Z%@�ZK@�Z ��Z
!�V� �Y� 
i � i� *i� :i� Ji � Zi� ji� zi�a�ioDEBU{�$v� u��;q��"F7O�50CAB��6��CV�z� 
fr����u kњw�!�w�!�w�1�w �1�w%A�wKA�w��p\0��"3LAB"2�|EwЄ�҂�3 ��*�SERV�EN� � $nq�_NAǁ!_�PO����` f�E�P�_MRA��� �d  T���EcRR����~ TYi���RI�V"0�S��TOQ�T)PL��T��Ѕ6 ����J � p�PTl X���_V1�b�Q���#��2�2+�����/@�8�p��5�$W��V�j��VN�[�$�@@�� �S���Q�	E�HELL_CFG�N� 5%�Bo_BAS��SRvp\0�K� �S��TJϐ1a�%Α2�U3�4�5�6�e7�8�RO࠘��� � NL:�3AqBn��АACKwv ��)�o��0u0iႩ7_PU2�COq��OU��P��ӕ������TP�_KcAR�0��REm��� P����QUE�٩��@���CST?OPI_ALzs���� �TĠ�� SE�M[�w�k�Mw�y�T�Y��SO`��DI����Є�=�װ_T}MK�MANRQζ� E��$KEYSWITCH���Ѱ��HE��BE�AT���EpLE(����&�U��Fd���|��SO_HOM� �O��REF�@PR�i��R� ��C@�O0�p ECO���� _IOCM�4M�k������'�O� �D�!ۧH�U��;�M�7��@�3FORC�ߣ�� ��OM>q � @Etx*k�U#Po1B�O��o3B�4x_�S�NPX_AS���; 0ݐADD��(��$SIZߡ$�VAR�TIPRr�q�G�A(ҷ��@
�˨r�t�50�SV��XC����FRIF��R��S%�7�x���N�FѲEАO� x6�PSIڂTEC*�.%CSGL=�T�"�0�&�V�D��>�ST�MT
�o�P\�ByW�@?�SHOWw���P�SV� K�w� ���A00�0 �Q��K���O���_���Ti���5��6��7��8��9��A����@6������20��F�� 
 ����U ����� �����0�� �J@��:�1�G�1T�1a�1n�1�{�1��2��2��2���2��2��2�2��2 �2-�2:�2�G�2T�2a�2n�2�{�2��3��3��3���3��3��3�3��3 �3-�3:�3�G�3T�3a�3n�3�{�3��454��4���4��4��4�4��4 �4-�4:�4�G�4T�4a�4n�4�{�4��555��5���5��5��5�5��5 �5-�5:�5�G�5T�5a�5n�5�{�5��656��6���6��6��6�6��6 �6-�6:�6�G�6T�6a�6n�6�{�6��757��7���7��7��7�7��7 �7-�7:�7�G�7T�7a�7n�7j{�7��
��VP$��UPD��  ��P���x�YSL}O��� � ��`հ�����QTAS�8sTƠ��ALU}U�����CU��WFdQIgD_Lѳ�UHI�Z�I�$FILE_�Σ�T�$u�_VS�A��� h��+`E_BLCK(�8bg�>AhD_CPUQi�� Qi���Sod_R1�ɢ�R ��
PWl,�d� �aLA��S���c�a�dRUN 5��a�d�a�d��5��a��d�a�d �T�pA�CC���X ;-$&qLEN~�3t���&p����Iѱ
�L�OW_AXI(�F)1&q�T2mwM��ɢ����I����Q�yGTOR.�&p�{DW�<�s�LACE���p&p�����_MAu�p�v�u�w�qTCV�|��wTڱ�;�1�<� �t?�_��s?�J�����M��ӠJ����u���u2q2�����ؾ��s�pJKцVK�~�か��3ՃJ0l���JJ�JJ��AAL�����e4�5Xr;�N1B�PN��	��tL�p_k�Ϊ��*!q���{ `5`GROU�P�Y�ӲB$�NFLI�C�ө�REQUI;REv�EBUV�"q���кp2���#pɖx!qxг�� \��/APPRՐC���p�
!�EN�CLOz�,�S_M ���A��u
!q��� 䆣�MC�r;�Xr|�_MGц�C��,`���N��p��BRK��N�OL������Rϰ_CLI��է����JޠѤP��p��p���p;��pD��p6�K���8��3��"q���G� ҒMr:ql�<Gqz�PATHv���@����Rx�������pCNR�CA��է�6��IN%rUC�pwQZ�Cd�UM�Yop�����QE:p�Gp������PAYLOA�ͧJ2LHPR_A	NqQ�L�`[�W�K��g���R_F2LS3HRё�LO\�������ACRL�_�����޷C�XrH��P"�$H���F�LEX�I!pJ>%u� :2Dv �p4�K�GYq�pPbt|F1Kљխ׃� ������E�� ��/�A�S�e�w��� ��y���ф���蘏��H��J�ÊT���X�� ��υ ��څ��[�� ��
�� �)��;�D��V�h�z�Y�J��� � �������QIPcAT��ё��EL4�S �ؘJ���ߐ;JE��CTRޱ���TN��F�ɗHA_ND_VBp��ܹP`�� $&�F20��K��ШRSW��X��j��� $$M��}�R��E��Uw�H��sA�PH����QD���A���P��A��AAɫ���j`��D���DɫP��G�`1)S�T��9!��9!N̨DY�`���|�Y�� ��KыǦ�J�ч�s�U�ХP��&�/�8��A�J�S�=��� �; �t�.R66N�/QA'SYM����Ґ�����Խ��ٿ_SH �����筈4��+�=�O�JV��h�'C�I����_VI��dHN�u@V_UNI�ÉD���J҅�B�% �B�̦D�ųD�F�̓�@�������*Uc�Ԓ�Շ��H�`���XQEN� v�D)IɠS�OwT Y�YPN��� ��I�1A��äQ�`Bc�S`�  p�a.a� � -ME����R4'R�1TkPPT�0) ���Qz�~���0�X�a	iT@� $DUMMY1���$PS_��RF��ЈP$Pf�aL�A��YP�jb�S?$GLB_T>mU��e�PpQ p���Q�c X	�ɗ`�ST���ߐSBR��M2�1_V��8$SV_ER��OÐ�c�cSCL�`�bA5�O�R�TPT O�P � 7D �`OB���LO˰&uq9c�`r��0�SYSqADqR�TP�PTCHb � ,&����oW_NA���t�z�9SR���l =��M�u` �ys�u~�s��s� ����������0� )�T�"�5�~���B�����s�?�?�?DY�XOSCRE)�p��ȐST[�s}��P!��tY�r _:� Aq� T	��` ob��a`�l��Ҥ��jg�c�O� IS��c��UY�UE�T�# �ñjp^`Sq��RSM_iqmUUNEXCEPlV֑XPS_�a����޳���8�޳R�COU�Ғ�S� 1�d�UE�tҘR�b9�PRO�GM� FL�$CU�`PO?Q�д��I_�PH�� �s 8џ�_HEP������PRY ?��`Ab_�?dGb���OUS�� � �@�`v$BUT�T�RV`��COL�UM��U3�SERyVx��PANE� �q��P@GEU��<�F���q)$H�ELPB�l2ETER��)_��m�Am� ��l���l�0l�0l�L0Q�INf��S@QN0�� ǧ1�����ޠ �)�LNNkr� ��`T�_B�μ�$H�b TE�X�*��ja>�RELV��DIP>�P�"�5M�M3�?,i�0�аN�jae���US�RVIEWq� �<�`�PU�PN�FI� ��FOCU�P��PRIa0mx@`(Q��TRIPzq�m�UNP�T�� f0��mUWAR�NlU��SRTOLJ�u���3�O�3wORN3�RAU�r6�TK�vw�VI͑~�U� $V��PATH��V�CA;CH�LOG�נ�LIM�B���xv���HOST�r�!�R��R<�OBOYT�s��IM�� gdS�P} 2����a���a���VCPU_AVgAILeb��EX��!W1N��=�>f1?e�1?e1 n�S����P$BACKL�AS��u�n���p��  fPC�3�@_$TOOL�t$n��_JMPd� �<���U$SS�C6���SHIF ��SރP`V��tĐG�R�+�P�OSUR�W�PRADI��P�_cb���|a�Qzr�|�LU�A$OUTPUT_BMc�J�IM���2��=@zr��TIL��SCOL��C����ҭ�� �����������o�Bod5�?��Ȧ2Ƣ��0�T���vyD�JU2��� �WA�ITU����n���%���NE>u�YBO�� �� �$UPvtfaSB�	T;PE/�NEC���@ �ؐ�`0�R6�@(�Q��� ش�SBL�TM[��q��9p����.p�OP��MA]Sf�_DO�rdATZpD�J����Zp>�DELAYng�JOذ��q�3�����v0��vx��,d9pY_���	�7"\��цr�P? �O�ZwABC�u� ���c"�ӛ�
N��$$�C��������!�PN�� � VIRqT���/� ABSf��u�1 �%�� < �!�/�/??0?B? T?f?x?�?�?�?�?�? �?�?OO,O>OPObO tO�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�_ oo $o6oHoZolo~o�o�o �o�o�o�o�o{� ���AXLMT�s���#  �tIN8&8qtPREO���+vupXuLARM�RECOV �)XrzujF ް%s   d�������7�I�[�m�~�, �
�/��vNG5� ��+	 =#��
ڏ�� PPLIMC5�?�%upՁ�Handl�ingTool �-� 
V7.7�0P/36 ���
]�_SW2�D�Fy0j�W� 43Y��J�9�K�7DA7�?����
&�X�e�	-�None���J����� �T7o�	�rP_��Viu�6s��UT�Oz"�,tTy.�HGAPON� %��!.��U��D 1�y� t�x�����y.��K�Q 1�{  THp������	��p�uq��"�"� �!��H�եw��HTTHKY��"ٯ���� u�����󿽿Ͽ��� ��)�;�M�_�qσ� ���Ϲ��������� %�7�I�[�m�ߑ��� �����������!�3� E�W�i�{������� ��������/�A�S� e�w������������� ��+=Oas ������� '9K]o�� ������/#/ 5/G/Y/k/}/�/�/�/ �/�/�/�/??1?C? U?g?y?�?�?�?�?�? �?�?	OO-O?OQOcO uO�O�O�O�O�O�O�Ƹ�TOĀ��DO?_CLEAND����{SNM  ɋ����_�_�_�_o��_DSPDRYR�_&��HI!��]@�_}o �o�o�o�o�o�o�o�1CU��MAX@ �bTQNQS�sqXbT�B�o�B���PLUG�Gb�cWo��PRC*4`B�P]klo^��rO�r=o��SEGF;�K�+�6��_�_�}�������ŏ�0�LAPZom�/��+�=� O�a�s���������͟�ߟ�6�TOTAL��v�y6�USENU
Z�g� HXL�NR���RG_STRIN�G 13�
��M,�S�
~��_ITEM1��  n󝬯��Я� ����*�<�N�`�r� ��������̿޿���I/O SI�GNAL��T�ryout Mo{de��InpB��Simulate�d��OutT��OVERRW` �= 100��I?n cyclHŕ��Prog Ab�or^Õ�>�St�atus��	Heartbeat���MH Faul<����Aler��� ��'�9�K�]�o߁��ߥ� ^S��^Q ��������,�>�P� b�t��������������(�:���WOR9���r���L����� ��������*< N`r�������PO���� ���9K]o�� ������/#/�5/G/Y/k/}/�/DEV� -�/�/�/ ??)?;?M?_?q?�? �?�?�?�?�?�?OO|%O7OPALT�� ^A��8O�O�O�O�O�O �O�O__(_:_L_^_�p_�_�_�_�_�_LOGRIxp��avO�_*o <oNo`oro�o�o�o�o �o�o�o&8J\n�_*�R�ݦqo ������(�:� L�^�p���������ʏ�܏� ���PREGbNK��$�r����� ����̟ޟ���&� 8�J�\�n���������~��$ARG_r��D ?	������� � 	$�	[�]���.���SBN_CONF�IG ��L��K�F�CII_S�AVE  ��k�b��TCELL�SETUP ���%  OME_�IO��%MO�V_H��¿ȿRE�P�|��UTOB�ACK��V�FRA:\8�� �8���'`��8�c�,�INI�a@8�^�,�MESSAGz�����|���ODE_D���}�C���O� ��,�P�AUS!��� ((O��J�\� F�|�jߠߎ��߲��� ������B�0�f�t��%�*TSK  �5ݒϕ�/�UPDT�����d����XS�CRDCFG 1v��� �������&�8�J�\�n� ��\�n���������� "��F��j|�����/e�2�G�ROUN����U�P_NAܰ��	�2��_ED��1�
��
 �%-BCKEDT-�0�}��pg�ӰQ-2�p8�/�/�8���g2���E/��/��/~/��ED3n/&/�/J/�\.�/"?�/�/ED4 ?�/?�/\.[?�?5?G?ED5�?n?#O�?�\.�?jO�?�?ED6 ZOO�O6O\.�O_}O�OED7�O�Ok_�O�\.G_�_!_3_ED8�_�o�]-�_Vo�_�_ED9Fo�_�o�"o]-�o�oio{oCRoY_Vh�]1��{� LNO_D�ELGE_U�NUSE	LA�L_OUT �V��WD_AB�OR���~�5�IT_R_RTN�ǀH�ONONS)Ю������CAM_PAR�AM 1����
� 8
SONY� XC-56 2�34567890�Y �f�@����?�W�( С���8�h�х�ڎ��HR5ǃ��	���R570�B�Affފ������ڟ� ǟ�"���F�X�3�|����i���į!�CE__RIA_I����5��F��;�Я� ���GP 1]����s�����V�C󠸾�����CO�C ��(���ǀC8��@��H̺�CCX����Ch꺰p��x���� +C�����Ⱥ���+�=�G��ށ��HE>/pONFIG=�f��G_PRI 1�B�$r�����������(�~�CHKoPAUS�� 1���� ,wuj�|ߎ� �߲����������� 0�B�T�f�x����D�O���T���_MORGRP �2?� �\�� 	 �,��P�>� t�b���5�����eҒ.�?a�a�����K(���d�P�V��a�-`�/A�

s��������b&�i��ܦP�DB�����)
�mc:cpmid�bg��:� � -�-y���p��U   ��  .s/3�� ��d�~���~��{C�e�*/��/��{g�+/���uf/s/i��u/�
DEF ̋(K�)�b buf.txt�/�/���_MC������d,53����|ʇ�Cz  B��p�B��FB�8��B��~C� �Cޢ�D3��u
q�Dzl'D�:�"DrBE�NNEA7E�V�ߓ=F�pg�F=C�F�e,�G���Gp��OG�/�	ބ	6:����4���U(D~���/�	�ʄ3@à1zTB��D�V@a  E�I�5� F*�� F�G$ˀF�[� GR�kNG�l��G��G���&H��G?֓�H��߃]���  >�33 ��ށ�  n4^��@߂5Y�Ed���A��=L��?<#�
 ���_�*2RSMOF�S��.^�9T1>��DE ��l� 
 Q�;�P � 0_*_>TES�T�"__��R�(��#o^6C@A�KY�B�Qo2I��B�0��� �C�qeT��pFPROG �%�S�o�gI�qR�u����dKEY_TOBL  6��y�� �	
��� !"#$%&'�()*+,-./�01��:;<=>�?@ABC� GH�IJKLMNOP�QRSTUVWX�YZ[\]^_`�abcdefgh�ijklmnop�qrstuvwx�yz{|}~�����������������������������������������������������������������������������q��͓���������������������������������耇����������������������Eъ`LCK��l���`�`STAT��c_AUTO_�DO��O�IN?DT_ENB;���1R�QY�K�T2�����STO�~��TR�L�`LETE��ފ_SCREEN� jkc�sc 	�UπMMENU 1i?  <�l�o l�K�u���FS���� 柽�ϟ���R�)� ;�a���q���Я���� �ݯ��N�%�7��� [�m�������ɿ�ٿ �8��!�n�E�W�}� �ύϟ�������"��� �1�j�A�Sߠ�w߉� �߭߿�������T� +�=��a�s����� �������>��'�M� ��]�o����������� ��:#p)+�_MANUALӏގ�DBCOu�RI�G�$�DBNUM�LIM�,1e
��PXWORK 1k�_-<_pN`r�TB_�  m��Y0�__AWAY��1�G�@b=�P�_A!L� =���YҀ��t`�_�  1!�[_ , 

:�&d2/o/�&�Mt�I�ZP�@P�#ONT�IM��d��&�
�e#MOT�NEND�o$RECORD 1'kqU2)?�!�O�?1 -?&k�k?}?�?�?88 �?�???�?c?O*O<O �?�?rO�?�OO�O�O �O�O�O_�O8_�O\_ n_�_�__�_%_�_I_ �_o"o4o�_Xo�_|o �_�o�o�o�oEo�oio �oBTfx�o� �/����� >�)�7�t�� pu��� ��-��͏ۏ����� N�`�Ϗ��o����)� ;������8���\� ˟ݟ����;�Q�گI� ��m��4�F�X���TOLERENC��B�	"�L���� CS_CFG �( +x'dM�C:\��L%04�d.CSVY� clֿx#A ��CH�z _/x.�G���},��RC_OUT )�- z/��?SGN *��"���#�19�-JUL-25 �13:08��27-MAY���4:3��]� Z�t�����x.�����pa�m��P�JP��k�VE�RSION ���V2.0.�11~+EFLOG�IC 1+� 	d��ٓ���p�PROG_ENqB�2��ULS�'� �p�_WRS�TJN� ��"�E�MO_OPT_S�L ?	�]�
 	R575x#V?�74D�6E�7E�#50i�d�o�2E�d���j�"�TO  �.����k�V_� E�X�d�% �PA�TH A��A�\��M�_�~+ICTZ�F�, '�>`�eg��}��STBF_TTS��(�	��Eм`����� MAU��ߧ"MKSW��- )��},t���.�!��]l� R�v������4SBL_FAU�Ly�/��#GP�MSK�ߧ"TDI�A��0����`����!1234567890xS�l�P�����// %/7/I/[/m//�/�/��/�/�/L0PV ���/� 2?X?j?|?�?�?�?�? �?�?�?OO0OBOTO8fO8<x�UMP$�I�3 �ATR>㜢O�@PME���OY�_TEMP��ÈÓ3��4��DUN�I	�w�YN_BR�K 1��x�EMGDI_STA	����_�LPNC2_S_CR 27[� �_�_�_�_�&�_�_o` o2or�nSUQ13y_ +?|o�o�o�olRTd47[�Q��o�o ���_>Pbt�� �������(� :�L�^�p������� ? Ǐُ�0�,p��+� =�O�a�s��������� ͟ߟ���'�9�K� ]�o���������ɯ� ����#�5�G�Y�k� }�������ſ׿��� ��1�C�U�g�yϋ� ��ׯ��������	�� -�?�Q�c�u߇ߙ߫� ����������)�;� M�_�q��ϧ���� ������%�7�I�[� m�������������� ��!3EW��{ ������� /ASew�� �����//+/ =/wa/s/�/�/�/�/ �/�/�/??'?9?K? ]?o?�?�?�?�?�?�? �?�?OK/5OGOYOkO }O�O�O�O�O�O�O�O __1_C_U_g_y_�_��_�_�gETMODoE 15'Efa t|�_Gg�RROR_PROoG %�Z%����HogTABLE  �[1O�o�o�o��ZRRSEV_N�UM �R  ���Q�`a_A�UTO_ENB � u�SZd_NON�a 6�[�Q�b_  *�6p�6p%�6p�6p�`+5pO8astHIS�cXa��P{_ALM 1]7�[ ���6|6`+t���&��8�J�x_�bp  ��[4q�R���PT�CP_VER �!�Z!6oZ�$EX�TLOG_REQ�v�y�SIZ��܄TOL  �XaDz�r�=#{�
ނ_BWDo�p%��fQ���_DI?�7 8'Et�TxXa b[�STEPg��y��P��OP_DO�v$v`FEAT?URE 9'EQ���QHan�dlingToo�l � DER �Englis�h Dictio�nary�7 (�RAA Vi�s"� Masteyr���
TE0��nalog I/yO��p1
0��uto Soft�ware Upd7ateb� "/�k��matic Ba�ckup
�d
�!��ground EditB��  25L�CameraT�F�X� "Lo��elylT��L, P��7omm9�shۡ�oh600��cou�Θ�uct��p�pa{ne� DIF����tyle seolectѡ- /��Con��9�oni�tor��Hd�t�r�Reliab�T�ϣ(R-D?iagnos��Q��	�H�Dual C�heck Safety UIFc��Enhanced� Rob Ser�v��q �v	�ԸUser Frܿ��T_i�xt�. DIO f�f�i�� )�\�en]dܰErru�L��O  prנ*�rO��� @���EN�FCTN Men�uİv����.fd�`�TP In?�f�aco�  
E�G���p;�k Exc�ذg�C��Hig�h-SpeܰSk}i��  Par+��H���mmuni�c��ons��\a�p��urf�?�X�t�\h8U���c�onnZ�2Т !��Incr��stqr)�8��M-6��KAREL Cmod. L��ua���}��B�Run-T]i�Env�(<Ш@�I�<�+��s��S�/W�"H�L?icense����� ad���ogBo�ok(Sy>�m)�	���"MAC�ROs,��/Of�fse\�f����H��!�Y�M1�Me�chStop P�rotZ�3� 5�
�Mi4�Shi�f\��B6S�M�ixܰQ����H�M�ode Swit�chY�Mok���.J�� ��Mt�Q�g��� �5��ulti�-T������)�Po=sj�Regi>����  ! �PA�t� Fun1��6isB/��R�NumⰈY�3�G�P/��� �Adju��	�/23HS�)� o(�8��tatu���AD� ��RDMޱot��scove&� �#e�v�㱗��uest 867.���o�\���SNPX� b��Y���)�Li�br%�
�rt ID���� "����.S��o� ��s in �VCCM������ j�����㣀/�I�� 710�TMILIBX����g�Acc����C{/2�TPTX�� �Teln��Y@�����K�PCUnexceptܰ/motn�� �������\m72�5����w�5���  �h640SP CSXC�i � j*��� RIN��We����50,��v9rl�زmen" ��fiP-�a���P���Grid{�pl?ay F O/���? ��ELR;�|�2�0��ORDK�s�ciiw�load��41d�st�Psatd��CycT��h���oriɰ:�7�c Data� qu6�2�0�*�����n��FRLamc�~K�HMI De��1(����k�PC�φ��Passwordn�644��Sp������D#YELLO�W BO�	?1�A;rc%�visu����#ti�Op�^�!k 2��aO�po��3 t��ֶT1o���f��HT��xy�^	�   $�t۠�ig��10Ơ 4�1\+�JPN A�RCPSU PR�+�8b!OL0S;up�2fil� �!p��E@-�;�croc��82��v���$ 1�2jSS0e4�t�ex-� I�7�Soz��tf�ssag�� e��У�P��,���� "Tc VirtȻ�v�!����dp�n�
�J3�SH�ADf0MOVE �T�MOS O �TԠget_�var failCs l�>PU~1E����� Hold B�us %�h��VI�S UPDATE� IRTORCH�MA A�{�vYWE�LDTV S ]�D~tS: R741���ouiPb}�y��B�ACKGROUND EDIT "R�C$REPTCD �CAN CRAS�H FRVR 6�2z1�SCra��s� 2-D��r )� "��$FNO �NOT RE��RwED �` m ���JO� QUIC�KaPOP FLE�N m41S�Loyc��gRTIMQ%�~#�FPLN: FG���pl m�r`�M�D DEVICE� ASSERT WIT PCV;P�B�AN#aACCE�SS M .pcv��Jo��Qui±��KbldmgUS�B$ ��t & r/emov�� Pg�SMB NUL� \;a|�FIX��C���ACHIN,QOL��`MO OPT �ՠa��PPOST<0�WDU C�wQ7Add�`ad���0kio�2��$P�`�W\0.$0`O�I�N&�P:fix �CPMO-046� issueC�J�/aO-�0�r130�Т- ��vRSET� VARIABL�ES-P{��R3D �m��view d2��M��&�ea���}b��of FD�5�P:N@x OS-91y0`�h sc���mt��s t�lo���7 WA�PZ�3 CNT0 T�/"�sImR�)�ca �P�u��POT:Wh�enapewB�ST�Y E�{1t��pt�KQdo GET_��p �p��VMGRw LOl�REAd0C~QW�~1�(�l�s�\gD�ECTpLp�ING IMPR�DR(p+PB�PRO�GRAM�ERIP�E:STARTU�� AIN-;�ӠM>/ASCIIzPÂ�OF Lq�DPT�TB: N�pML�$me P���`:vx�mo&�allW`\!�ӤTorc�A��U�HC�iLpԸth:�`n�@ ch��/8GEA�!�tou͐��RCal��k�Si�gn`� ND�ԗT�hresh123�`��09p : M�SG_P�+0er�  �Q�Aܠze�ron��0 H8�5��RImA�n�2�D��rc�0I��O3MEa`�pONaP5��  נSREG:�FF-Д� ]�'���K�ANJI��n��Jr��c�0asn d�!�OA immc �I�NISITALI�ZATI����~1w�em����dr+� �LB A�UWqmiwnim�rec[��c!�R���m$�ro� -1>ѮS�ܰi�r��@ұJ�1pdETw⌀ 5`?�I�ow �u��< se 1lc��YbPM���p�Q`���R`vR&�lu\�3�Re 0�4q�q�1#���m <a�a�rn��ঁBox� fo��*PRWR�I�PW�S��v�09� F�pup�de/-rel2 d�p� �j��`━betw=e��IND Q����igE snap�|�us��spo wTME��TPD#��DO�p#aHANDL 1\k�`vR��
ȀD�ny�S�v�Y�operabil8� �T*�: H � 	l\p��Vq�b�R�< �p�a*�c&2O�`F�A,�.�-QV7. �f.v��GT�p�i�s��� ɠtm�Line-Re�mark �� R�M-�` W�#SPA�TH SA+PLO?OS UIFc�+5�f fig�pGLA�����Vrp������U��0ther�V� OTrac���tW�\b�s7��d�t��� n�@  ���3:����dK�y��its k8�d�PayR!�[2]�ü1: ug��s��dow�XQ��0IS�q�qE�MCHK EXC�E C���MF �+�Xah�� 35C\k��)���QBt�@���'b���[�c����e �`k�S�� GBUGr��cD$`�PETp���f�c�4��0XPANSIN��DIG��@OoP�metTCCRG �EN��CEMENiT�A M̀K {���`H GUNCHsG �`� EXT�Ph�2�bQS�93 �wP8�x�ORYLE{AKq  H5g�yq�PLC WRD7N R �O /u�Q�SPE=p��G*�V� ��$�tn720]\3pGRI��A��rT�PMC ET�H��pSU7p�` � j5/n�PEN�S�PN,��*P o{nt�`BROW�`�!sRMV ADDfz CN qDC��~�PT3 ALA2@� ���pSVGN EARLY�R��Ű�H57�GaJL�AYҀE (@M��PPD�p*@H�S� I`P�OUCH�8���V�F�q�co�mH�x ��ERRO=R� DE nJ��{RO�CURS�8pI��N4q�-�158n7�RSR	 xP#aUp���Rq
y�T�Fz�;�pk���t�� gՂ�B��SY RUNN��  a�`�BR7KCT�!RO�p3@� \apSТ�AXxP���h8+ q��ISSUr} sPX��PTSI�K1M�10_�IPSAF�ETY Ck�ECK[��Á������p<#X�� �TWD2��@�@�INV��D' ZOp�5X���t�DUALy� "�M6�0�"rF#�E���dPdNDEX� F�t*UF��"Pʀ�0sFRV�O117 A�PT�6�KtqFALPT�P2477D6_�Pܞ!;HIG� CC��t;SNPX� MAM��tq�d~�Vq�q#�
"��DET�EC�Tq*@RRU@�qA�P�5p�9 y�!)<9���7T��P?ds� k�	𐱬!Q���� t\�4A�;A0�2 "Ke@" 8@HI�qXF8@|4@H�PRDC"�
�aMB8@�IXF�b� ��zOX@8@���a�G}E<�B�Ccscr�J8@��Ndctrld. �A�NZE�A5��Q���!�`�Df8@�`m�8�78�Q-;� ���� rm`�
��PR6̠78�@RI8@0q�Q (~\Mp��0t��!{B8@\tQ<OX*�St0�3hB3nO�Vstp�A�@LCF�L���� �Rplcf����J8@�WTamai0�E8@mubov2_mi TA�O�S8@U`T[tT�A�qPr674xSShape Gen��8@j�I�[R�`�@8@1T����%q (u8@��II�^�Q~C�a�[X8@;Ynrsg0�4� g� 4�CtMr68@��r5hB5�zVnre[tsp "r�Po��wng0bGCRE�Ka�ޠ�DAT��E�k�creat.�q�M�a�oksqgtpad1P��(�tputZj�{�������܆28@����Q̢���sl�o��� �hexH�TB�8�ď�keyH�8@�#pmZb�NR�u7A+�nrgc8@UQ�pp�b�UZ�dp0aj921�xSpl.Coll أcq�\A��RNq�UfA� (J�8@ip�_@�WA��_�Y��a7hB�7�ͦtp[� "�TCLS9oKb��cGlskyh[��s�pkckZd���$�TQ`���dA�rx�710a�- KAREL �Use Sp�F'CTN9�a�7l�0s0a�� (���a��~C�8@��MI��c8hB8�"   �8@ �v	�v	�   lmatea99�qM�����E�mcclm5�C�LM;�� �j��E�et���aLM	�h�ya�sp,���mc_mot�B�N��8@H����Q��su'��Q�ȕ�8䅮���joi#��<���A_log�Z����trc�B����ve�ϓ�v��QWX��6��finderxSCenter F1�lSw520��ha6r6X� (<�r,�Q�Ձfi�Q �NH0�I��ۡ���A8@uL��tq~�a "FNDRV������etguid�UID�C8@����������TA@�nuf�;��P���ƞC�B��_z�Ӡo��qG����x��l���fndrTY8��2䁴tcp"�,qOCP MF�}38@g517��6s38� E��gf6��(��K���Q��-�X��A�tm6�P�İ��Q����	�͘��tm�Ĵ�b8@ej��TAiex��aP�Aa����cprm�A��>l�_vars��
 ��dwc7 TS��/�6恴ma7AF�Gro�up| sk ExchangJ 8@�VMASK H5�0�H593 H0aHi5@� 6� 58�!�9�!8\�!4�!2���"(�/��;OMI(� `@a0hB0�ՁU4U1#SK(x2�Q$�0I�h��)�mq��bWzR�Displ/ayImQ@vJ40j�Q8aJ�!(P���;� 0a��0���� 40;�qvl "�DQVL�D쌞�q vBXa`�uGHq�OsC��avrdq�O�xE�sim�K40sJst]��uDdX@TRgOyB�Bv40)�wA~���E��Easy Nor�mal Util�(in�K�11 J553m�0b2v�Q(lV40xU)���������k986#8�Uϕ�|�rP "NO�R��dw d.a}oKksu�O�W���OY�W`�j�0�6�H� menu�uyP6�M�`wRX�Rw577V�90 �RoJ989}�49bt\�`(�fity������e�<?��Vsm	h`��8��C0�Sv��q�8���w�pn? "MHMN<��� �x�Ay`�o�3�u�`f�І�x�t��tRzQ�0�LV��vP�tm���|"I�1{oPx �2|����I�3I/B�odst�Ǐًmn����}e�nsu_�L<���h�!!��Rt��hus�erp��0Ҹ�ʐc M�_l�xP�oe��рp�oper����xdetbo/�l>�x�� �Ps$p�`���OPy?dspweb͓���z'R��u�Rr10!1&S՟{t�`2�Z�4�30������`4�
�4�5��KQ�m[T��dUCalG40` �Q)p40}�����9;���DA�� sv	LATAumpd�\bbk968��68c�fbl�41969y�9�|�D����bd� "BBOX�êM��schedx����m�setuM:�����ff���40���n�41�ϒ�40q�ccol��|�1�xc������li��X�0����j��&�8�4 <�ro5�TP E�#��ryK42r��;�s(T+Q �Rec'� ʈ1Iw�84�����ޠAk971��71��;���parecjo��QNS�[T����dXrail| n�agek�M ,QT2 *� (�ĜR%<x�80!bh��p��4��4�yDgl��paxrmr "�XRM�g�l�brf{���n��kl��9?turbsp���8��- �l015	�g�625C�Mh�+π��)89��	+��B6@��o�ҹ��x�7�q�40����pd "�TSPD�=��tsgl��l�:dQ���8Bct���K�vrE�aܮ����~�  �!����21�`( �AAVM �2�0� �@fd TUP� him (J545 l)�`�8 616 %��VCAM ���CLIO (�0u:�5&  (F\ OMSC �Rt"PBs?STYL�D!�28 :2\ NRE� F2h SCH6p�DCSU t�psh ORgSR �rD!04�S�EIOC& \�fxh 542 L�EX"� ESET�n�8!H ��sh8 7�H �MASK��Ø"7>��OCO*`x�!03"6�!/4�00:66$ G639�.6[8LCH!6OP�LGR703
5MHCR��0C� (! ڢ06�A.f8!54�
��00DSWb 5�88�180 �h!37� 88 (D�"0�2C24���27 q�9�25��2-6�05���9PRST� bBFRDM�ES�!zB�930� _ NBA  �6� HLB 3 �(~!SM�@ Co}n� SPVC ��8!20z��TCP� aram\�TMIL A��@P�ACETPTX ��@p TELN �96��29�%UE�CK��r UFR�M et�P!OR� ORP IPL%C�SXC�0j�1CV�VF l FQH?TTP stA")�I#� CGHP8ZIGUI�0�hP�PGS Tool6� H8�@djZ��!�@�h!63�%�@3�2Q\�31 B�h!9�6�%R651�Rs��!53 TFADf�R41�8"1 ��oo�"9��417�75�"/@�P�VCT�O�@�U�!sh!80��%PRXY�R�!7�70 �b8 885' ol3P� L� а�di� �`ڳh LCxP{Q� TSS �b��26:����@CPEu �HT@VRC�~�tQNL ��@0�02 %��b	0dis� �`7 <��a\0l�T�`1 �`en�b�4 652�`)FU�02Q0Πo`p�PtLu�r4 $r5N�v�RU0p@nse�Q~Jp1 APFI[ �Jp3�g34�g40� alxrE1t4m4w46� ts �U0  7v�0O��r5��e�p7 p "sMw�a61:��r4��r5 QpwGr`�$��p8R�"sP`tQ�b�36w77�w8`�v83���r8�&:��p�Oq8�8 "rkeey8�9F��a90�91 p�#@��� �D�095�g97*pur�A1@d���P|PR�q1�0QplSq1p�#4��]a!s1@sl�༂8�Ӽ�\1�d1D�`��v�@{�14p:�ae��5 h2��`R�6ޣ��7�f1p@���d�YpCqd�ـd�1B�`uq��� Cu1< hOq� ��7ReU1$ ��u1�Pϱ� ��@-� WQ158 aose C��9 B>��60 82ń�p����4 (Wai ��`吢!��7E��m8�EU1P`ro9�<�1��<�2��<�	0 ��T��l�5J�l���cC���9%�MCR��P�2�`�Q�2@967�Q��8��9Z�2TPB��4�P�2P7U5@ࡈo���
�5�`U���3 w���?A�E�1��	c�qAwl��A�1>��512 f��1"�u5Р���a5p$B��56�+a��Q5h��Ұ�1 @��pp�b[�538 xaBP��|p�4�2�11/q�5�p�4U5�P16 (߲�Pz��0���8�P�����p�e5�`�e5(�/�P`bbAf>�X��$Z�U�5d��\� X�7 �	  ��8 kw_kv��79 ns�82 &�H5�� E6���p����h���È����3J"�`��4[ 3Ȥ59ѧ6�0)t���8��6D0$�.$�4 7��!����<�j670\tchk<�Ps��<�B<�90��7�<���<�	\K�<�q�Ӻ�A�C@<���q�<���<�t�ӛsg<�lc���FA<�H��<���<Я���<�hk��<Щ�B <е�o�<���<��K�<�dflr��<Ш��� ��o�`���D�;�<�gEvam�� ��B<г�oќ���<����KЀ�creex l����P��<���|�֭�j6<�s��prs.`���\���<�7�������fsgn0��P�b�t�at���<�L��1B !�sv�sch/  �Ser�vo S��ule�>�SVS��44`�1u�_<��� (��^��ched��,��0~��A\�� �� B����B�qA����cVj�� � 5�1<����Ә�p�css "ACS<�&(��6� �����c e�l���Q����to�rchms�<�- T�Ma`Ѵ���0�9 J5;598_ J681s�7� 8��b��<Чa����te,s�����p/�E�� m���ARC.�� 1�q�4�!=��C�tc��pA�@t���f� �F����7#�2x�S�E�r���UtmS�0960'���RC������� p��96G= '��"H5W����L���\f�� �PATb���`!4U�#!Stmt�E ��� �pMA�!p��8z�2?�in_<�X�(�r�X e/cW�����V����etd�l�vߏ\ovet�o���܏��mmonitr�\��|#F�0st��?.6a�`�PP���! Q8�!y`�`ame �Agrol�c�43��0 �p���01�� 25�  ��<� v	��v	�A@�818\n; <s�I�B�2>�pMPTP"��C>�1mocol��,� �CT�v�'!� �A����8P53��y`Touchs�s�`��<��J5���Ѩ`mP����n[PQ�a,�E��a��IP&
�Pth��A<�KF#R�m;�Qe�tth�THSR�'�q-�Rt��o "PGIO�#!$s�IS;wka�"WK��!v�MHqH54��%5w5n/�Sm/��B@ 7�*�da��8`!pw/Ac��tsnf Tk�/�#gb�a��u`��^m�`u��Zӭ�ܱQp�є�#���Ka$<��M��t5Qt Z�a<��dFS5GK����G�1or��dW��64��tPx���P ����x,��?$����P<�Z4e7�g "�SVGN.ox�co?py "CO;�Wj�$�O�A�9� "FS�G�ѧ�%7��_��f� wQSWF*!"(�sgatuɀ���_�
��tp_TPD4o��9�79�#d�p�?���h�GAT����!#��   �Гf�` ��"/� �w�Z� �b?6?� ����р ���E ���M� �c�hrT� �K6K� �s�ms� �o6�ѐ�gtdmen?3 �?���| ���mkpdtd2` ���, ���pdQ��X� ����� ���mvbkup. �[�C�<С��mkuno��sprp���mkl �44��s �niU��֞ �ldvrw���glg�4�� ��棑�n�aut7�.pб��旐 �ַ������su3� �Ǜ� �Ƿ�d ���\ �6�b2XՀ ��&�� �����A4�  ��B   946" ��fB�� �t\paic\?p4k947 ����F#���� �icta�s���pa`���c�c:�<��o�����g�en�� � ��F�l�np � ����stf@��1��wbO�c���p��`��߄�vri�� ��а�-T� ���p��flow� OPA�c��ow���R5�0qtS �#T� (A��4�#���pѣV�cu3�QF� ��SI�3ac����46����s&��pa��!!���� ���55�b �o�)�p���0娿
�af'cal3�P� ��f�P��}���`�f��m	�@��p�d�m�/���a/����$C`ѷ�� �! track\P� 0��ine/Rail� Tr�]TJ�69W�T  (L��8( `љT.�`�%��D��P�0� (��8�48 ��_ɛ�⇒4����(�� �3�b3���falV@ �NTf�0��%��Iin]0m���aen�������&?5�c@Itst3@��$���� `�,R9�%���0氱�%��popene�rs-OW dDev��F�M�6W���`|A�Pc"�l!esv�  �,��R��V$�Q���U�<�V$ �k9j �6�# �����%pa;op/!OPNU�8V ��2celL���8g_��/�6��tscG��$��V!�3�= 5vrop�ߡ�7`�n(`�V"2D��a V'O$:S9��� PumpE��jQ�@@�" ��!
��@бMSC #�@��)P��AC�`�<�� � v����� \mhplugB�@g�"7P��uK",)㠱io7�CJ0��\E�LIO q1g M7A93շ�5 q�9 t����4rb S�T��R��CPJ9899�P�LSE�' ��e C3Q(P �/O�v���o�P� ? 0I1�R���55��f�|I1`�tcmio���MIO�����Utc>o1"CL01V �YcBK`io��uM?���Sl�I0�ߢ�Eg" �o���f �tI4\onfdtI���e%�<p27�Inte�TB� CoMoo1E�R��(do554 (;r>Ex,��nR�##ipc�/>��qp	5���
oQé�1�pD����7/o���ra�pd�CDV_��rP�p֮��qp2cnd��s �p��a�o�r`� ��S��"�c�a�c�Ƃ�2kIԿ?A�pcCrt���or0�qd# ��"���3p+���D��<Џ��vr2k�0����AG�.+��cho�;�uC��(� �uV630�fwe Pmී�@���`��T�X�� ��d�chpC "_��(	�3������8����\p3��v����ш�9�3�1` �����low�[ͧ���chk���コ�s��s?Ө0�i�1 h���2��i�w����s?1*�-	�:�O��vr������0�'����PFRAPWat?1rneE�P�sp��& ac5� _A�rbo#�,�a��g� ������Qs<�ICSP+ 9_���<�� ��F�An9PH51IQ93 	7��HX6hQ]PVR`S5��fPR6 iQW�PR� (P!am S�u�"�A�I0�tpprg�0����`h�@2atk93�2�!��E�^��asc� "8�C��S>i�atp�"�d�@1I�
�g�dsblfl�tJA�QsableO Fau�P{C!���EV0ex/!DSB' (DC��t�$� p��X 7� �� 5��Q�t3*�~���td9� "!%�(5䆠�sb9኏���\�	�6#���@5�p$D@5�50-Adjust PointO"tVJ�Rs�z�䐄��!ȵX_�Yj��0\�sg��4��}7y�\�ada�"ADJ����j�Qetsh=a<�SHAP�sŭ'jpo�r4�t�!���$ ��C|�	Tkr!bRPKAR/Q�iagnosti�̀!O!vV66 JP`ew0�(�L����/�&krlde � ��PP���hU b�В�r3�Pp?q��D'BG2C��� �X �o�1U�� ��WXT`�@ipJCM�a�ipper Op�v`1Se}78 (MH GF� ;": �&##�� a�x�֕$��388C�����#
��9.�9C��g##PP	k�Q��8�!�_"$�" ��=0%�P��A $��_��#%0AQ�C~2 Mat.HandlE��!= &�pq MPL!GET�0�1(�3�T t&P�Sٰ'�B�1��B 0����&p��H��PP  �'p��@�C7PP	��TG�tD5�}m�q�Af�hnd "F_R � �����PP	   xT?Q���P7(Pa��To��(���?�pmpaO�˼JP ak925��2�`@O�JRpsQ`B2p�unLHP�Tgse��GSo1�O�W�QT`��v !�R�Ptp~�<��JRdmon.�@�̔V�!ns�hYvr �QJ�g�Q�o�jY�HS�~7sl�f ��pen�PDnR(R&���ɐ823'��ٔq�� �g� ���� 1�� S��: ? �c\sltQ�! |QE�P��a�rtPg��P�� �v��"SED�G8�s0�qtdgY T����vP` ho�s`<`����qc�`g
�e` o�w�a@oN"�ile6�H�e�e ̏nR�� �e! j517�>Ճ���J%��e�`��Q4��Q&�L�!F�J��=�o�5�z/l17@���_�œ��`C0C�?  ���LANG j��A��������gad���#�jp�.��4�Ē�ib���s�Ƒ�pa���&���j�539.f�,R�u� Env
 ������3H�z�J9�����h�Ф
�(����2�2�씤� (KL�n-T�imФ�⠤��p�3p�TS����\kl�UTIL"o���x�?r "QMGl��!p������1 "��S�T3�\kcm�no��SФT2���u�t�.�lreadc�}�exY�ܤ�r��E\��l��Фw�3��2C�*� -�C�D�@E!Ĥ� .��C� R cCV̴�Ҁ�\p��蠤��p�tbo�x��.�@�cycs�L�:�RBTE�ve�riOPTN E���;ӕ�k�e�ߦۘa�ߦ�hg�ߥ�D{PN��gp.v�|�r�ptlit���0�4��te\c�y����tmn�u3`�r���5UPDT����p���駣��ite >�� swto�,���oolB�F"��Y���Q��(q��gr�3��䪒��"�䴁w ������߳��s���@����������lS���bx "O�� ����l����P���A�l\t�� ������\��	�Col�e!��R C��r��&r� �m;`��Chan�g�Lq�T1 �rcAm3�"��
� 6���"����sP7���"�&�222��2dD457�<� CCFM�H�>�accda��Q�c' ��KÕ0���K!����mo!���,$ Á��!"
����/ �/����	Y�,$��)��,$sk����m rC%tS1,$+��k1�%unc.,$oñ�1��sub������1��cce�5/!&�� -/?-W/i&vs�}/ �%#�#�/�.C��/� C%
�@? U �&+��F�:qt�
pDЃ= D	  U�:�7�Dxmov.��P��DPvc5Q�tf�r@PeC_UYgeogbdtg_y[tu����P���PTUt�P�Sx�_�^z�_�\var��_�\xy�_�[pc�l`c�P���P�Ue~�Pgripsuao�skuti���ovfinfpo}��o�j�b!�P���Qud\�aX�P�Pc�\Rrp�Qnƅ�P�v�P)tm#qƆ�P�v�a+rog�a��\Q8�?a+rpal?a{�{spa���P�u�Q�tĊ_TZp�0�osipk�ag3r�ovlcl�ay(�:�t�pT�d �pu?a�c�A����@��KtKa�P����qT�f|rdm��{rin#r���s� �2�ě�|s�Pd�v�tvĈ�v�h�0��ystQn* џ�yt'�1�p���D�p�uϑ#�ul��@o�W6�2�siucpdl�]�o�vr�on��`1L�z�`\�r�΄�il3$|l4��ǉ#q54FyB�Տpg{�`���{wcmס<���wxfer�UY?tlk2pp߿UY�conv��sicn1v�Qʯxag��HώZ�lct`ao�=�p<��׭nit0믁��3������  ��� v	��v	$��alϑpm�r&�B�eWa��� f�%������I��� ��u�ͬ�KamT�f�0��c��w��roǁ#� 5�����?� sm�� y�a��y넑������ `����͐ϑ��p��m�Wa�1���A� 6�S�e�X��ψ�\Q}� ����������ĥw߉� 西߭���߮�#q0� �rs�ew���1�a��z긱n@�.�۲;��d������  }� Ad	T~$�1 p! P쥰e �e 	tlf@C�@�s/�  ?�����8� �x������reg.�C�=��o99 �~@����$F�EAT_INDE�X  z ���e� I�LECOMP �:���1!�!z$#SET�UP2 ;1%�;"�  N �f!$#_AP2BC�K 1<1) � �)��/�/  %�/�/e4 �/�/ >%�/$?�/H?�/U?~? ?�?1?�?�?g?�?�?  O2O�?VO�?zO�OO �O?O�OcO�O
_�O._ �OR_d_�O�__�_�_ M_�_q_oo�_<o�_ `o�_mo�o%o�oIo�o �oo�o8J�on �o��3�W�{ �"��F��j�|�� ��/�ď֏e������ 0���T��x������ =�ҟa������,��� P�b�񟆯�����K� �o�����:�ɯ^� ����#���G�ܿ� }�ϡ�6�H�׿l���@��ϝ���@)t Px/� 2� *.V1R��߅�*�@�`��F�j�T��PCr�|�߅�FR6:��"��V���z�T � !���K� ��q�SƏ*.Fߢ��	��Ӑ���^����STM ��'����S���iPen�dant PanelS���HI���9����U�������GIF 0;��������JPG��;��]�oR�
ARGN?AME.DTy�E>�\"���R�c	PANEL1Y�%>��e�w��2�A/�//���/�3_/�/� �/p/�/?�4�/I?��7?�/?�?TP�EINS.XML��?>:\�?t?�1C�ustom To�olbar�?Q��PASSWORD�g?w�FRS:\�:O�? %Pas�sword Config{OR��OSO �O�O��_�OB_T_�O x__�_�_=_�_a_�_ �_�_,o�_Po�_Io�o o�o9o�o�ooo�o (:�o^�o�# �G�k���6� �Z�l�������Ə U��y������D�ӏ h���a���-�Q�� �������@�R��v� ���)�;�Я_����� �*���N�ݯr���� ��7�̿޿m�ϑ�&� ��ǿ\�뿀��y϶� E���i���ߟ�4��� X�j��ώ�߲�A�S� ��w����B���f� �ߊ��+���O����� �����>�����t�� ��'�����]����� (��L��p�� 5�Yk �$� Z�~��C �g�/�2/�V/ ���//�/?/�/�/ u/
?�/.?@?�/d?�/ �?�?)?�?M?�?q?�? O�?<O�?5OrOO�O %O�O�O[O�OO_&_ �OJ_�On_�O_�_3_ �_W_�_�_�_"o�_Fo�Xo�_|oo�o�o�`��$FILE_DG�BCK 1<����`��� ( �)
S�UMMARY.DyG�oblMD:�o�*n`Diag� Summary�+8j
CONSLOG qn�=q�ConsoleO log�7kp�MEMCHECKФ�2��qMe�mory Dat�a3�;g� {)>�HADOW(������C�Shad�ow Chang�es���c-��)	FTP������=��qmmen�t TBD;�;g0�<�)ETHERNET0�`n�q~����=qEther�net �pfiguration���B`%�DCSVRF�/��'�@�C�%�� verify� allC��c1p{� �DIFF8�p�0�ůD�%Z�diffǯ{��q��1������J� �X�q�|�	�CH�GD�&�8�ͿD�ܯ�����2Ŀ�����R� `�yτ�GAD�.�@���D�����FY3�ϳ��ώZ� hρߌ�GAD$�6�H���D������UPDAT�ES.$�
�ckFORS:\"�c�>q�Updates �Listc�`{PS�RBWLD.CM���blN��e��pP�S_ROBOWEL\�6o+�=�loa��o ����&���J���n��� ��9��Jo��� "��X�|# �G�k�d�0 �T���/�C/ U/�y//�/�/>/�/ b/�/�/�/-?�/Q?�/ b?�??�?:?�?�?p? O�?)O;O�?_O�?�O O|O�OHO�OlO�O_ �O7_�O[_m_�O�_ _ �_�_V_�_z_o�_o Eo�_io�_zo�o.o�o Ro�o�o�o�oAS �ow�*��` ���+��O��s� �����8�͏ߏn�� ��'��� �]�쏁�� ����F�۟j������ 5�ğY�k�������� B����x�����C��үg�v��$FIL�E_N�PR]����Y�������MDONL�Y 1<��U� 
 ��ۿ(��� L��5���Y��}Ϗ� ϳ�B�����x�ߜ� 1�C���g��ϋ�ߘ� ��P���t�	���?� ��c�u���(���� ^�������$�M��� q� �����6���Z��� ��%��I[����2����VI�SBCK����ų�*.VD�*� OFR:\V� �Vision VD fileV d������� 	/./�R/�v/�// �/;/�/_/q/?�/*? <?�/`?�/�??�?�? I?�?m?OO�?8O�? \O�?�?�O!O�O�O�O �O{O_�O!_F_�Oj_ �O�_�_/_�_S_�_w_��_o~�MR_GR�P 1=��L~eC4  B�`�	 ��lo~li`�۬B��D���fnӺ�MT� ��� ����e`i`a�o�k hb�h�o�dcic.�N���L�/�K�.!M��M�H>a�E���|�i`@4���B��Az��?�Bf���9�f�l}A��U�A��A���lA�=A����p�l}F@� �qhq�y�~g�f�F6�D�Mq�D�� BT��/@���l}?pD�ޒ6���l����5��5����|�l}B���B��C�B�jZB�j�ZB}x�B�X�~e9�B��B(��A��}jA��cB��dl叐�A�����A�܏e�P����t�  @����@h0?�\	@�B������Ο ��+��O�:�_���`p�����eBH`� �ā��A`C0O���'�d
���Z��WZ�l�0/�FX
�A@����@�33@����\��[���ѿ�z ��񿋯�*��N�9��r�]ϖρ�<�G��=�<�m]�<�+=~�m�<c^��8e�N7��7ѷ7�x7;��51���	ߤ��?ߪ�d2^`Yb`�b`�J����F�`Үb`� b`�0�����C�^o�߂o�o�߸o ��o�� ]�(߁�l� ������������#� �G�2�k�V�{����� ����������1  ��-�)�� �����0T ?xc����� ��/')�'/M/_/ q/8��/�//�/�/�/ �/?#?
?G?2?k?V? �?z?�?�?�?�?�?O �?1OOUO@ORO�OvO �O�O�O�O��_��J� ���`_*�_N�_�O �_�_�_�_oo'oMo 8oqo\o�o�o�o�o�o �o�o�o7"[F jh�x�t� �!��E�0�B�{�f� ����Ï���ҏ��� �A�,�e�,/������ ���/�J����=� $�a�H�Z��������� ߯ʯ���9�$�]� H���l�����ɿ��ƿ ���#��O�OV� _z� D_V_��z_�Ϟ_�� �
�C�.�g�Rߋ�v� ���߬�����	���-� �Q�<�N��r��� ������)��M� 8�q�\����������� ������7"[F k�|�|���� ֟3�WBg� t�����/� ///S/>/w/b/�/�/ �/�/�/�/�/??=? (?:?s?:�LϦ?p��? �Ϧ� O��$O��T?]O HOZO�O~O�O�O�O�O �O�O_5_ _Y_D_}_ h_�_�_�_�_�_�_�_ o��@o
�go*owo�o �o�o�o�o�o	�o- *cN�r�� �����)�;�M� ��������ˏݏ ď��%��I�4�F� �j�����ǟ���֟ ��!��E�0�i�T��� x���ï�?�?��O� �?OO�t�>O���� ��ѿ��ο��+�� O�:�s�^σϩϔ��� ������� �9�$�6� o�6o��Zo��R����� �����5� �Y�D�}� h������������ �
�C�U��y����� d�����:����� +Q8u`��� ����;& _Jo����� �//گ4/��x�j/ 4��/X�n/|��/��/ �/!??E?0?B?{?f? �?�?�?�?�?�?�?O OAO,OeOPO�OtO�O �O���O�O_�O+__ O_:___�_p_�_�_�_ �_�_�_o ooKo6o ooZo�oZ��o�o�o�o ��xo
G2kR �������� �1��.�g�R���v� ����ӏ���	��-� �Q�/*/��N/��r/ �/ޟ�/��/)�D�M� 8�q�\����������� �گ���7�"�[�F� k���|�����ٿĿ�� �O�O�O��W�B�{�f� �ϊ��Ϯ�������� �A�,�e�P߉�t߆� �ߪ��ߪo��+�=� a��߅�p���� ������� �9�$�]� H���l����������� ����#G2W}�h�p��$FNO ������
F�0� �  #�1 �D|�� RM_�CHKTYP  �� �q�� ��� ��OM� _MsIN� m�����  X� SS�B_CFG >�� �~�Jl�Aj|�T�P_DEF_OW�  m���I�RCOM� ��$�GENOVRD_�DO����T[HR d�d�o_ENB� ��RAVC_GRP� 1?3� X �e/��/�/�/�/�/ �/�/�/? ?=?$?6? s?Z?�?~?�?�?�?�? �?O'OOKO2OoO�O hO�O�O�O�O�O�O��ROU? E� �q������8�?#�O__K_�m_o_ꐖ  D3A���_E�_q�@A��\Bȡ��R��>Y_�6 SMT<#FC-�Ufoxo�o�HOS�TC,1GY?[��_ 	�h�k��o�f�oyeCUgy�z1�������p	�anonymous�5�G�Y�k�w��o �o�o������ *�<��`�r������� ˏ	�����&�8� �������������ȯ گ���M��4�F�X� j�����ݟ��Ŀֿ� ��I�[�m�ρ�fϵ� �ϜϮ�����}���� �,�O�Pߟ�t߆ߘ� �߼���/�A�C�(� w�L�^�p����ϸ� ���������a�6�H� Z�l�~��������� ��9� 2DV�� z������#�� 
.@�������� �������// g</N/`/r/�/�� ��/�/�/?Qcu ��/[?��?�?�?�? �?)/�?O"O4OFOi? �/�/�O�O�O�O9m�a�ENT 1H[� P!^O_  `_?_._c_&_�_ J_�_n_�_�_�_o�_ )o�_Mooqo4o�oXo jo�o�o�o�o�o7 �om0�T�x �����3��W� �{�>���b���Տ�� �������A��e�(��:���^�����㟦�?QUICC0�̟ޟ?��1@��.�����2��l�~�߯!?ROUTER௼��ί/�!PCJO�G0��!19�2.168.0.�10	��GNAME� !�J!RO�BOT���NS_C�FG 1G�I ��Aut�o-starte�d/4FTP:? �Q?SOBχ?f�xϊ� �Ϯ��?�������+� ߿�P�b�t߆ߘ�6 �����(�J� �1� C�U�g�6ߋ����� ����x�	��-�?�Q� c� ?2?D?������� ��)��M_q ����:��� %t�����m�� ��������!/ 3/E/W/z{//�/�/ �/�/�/6HZ ?n/ S?�w?�?�?�?�?�/ �?�?OO<?=O�?aO sO�O�O�O�/
??.? 0O_d?9_K_]_o_�_ PO�_�_�_�_�O�_�_ #o5oGoYoko�O�O�O �O�_�o&_�o1 Cogy����o T��	��-�|o�o �o�o����o��Ϗ� ���)�;�M�_�q� �������˟ݟ�ÿ�T_ERR I������PDUSI�Z  �^����$�>=�WRD �?޵w��  �guest +�}�������ůׯ���SCD_GROU�P 2J� ��`�1��!��L9_���  ��>!�	 i-	�E���Q�E E�ATSWILIB�k�+��ST �4�@��1���L�FRS:аT�TP_AUTH �1K�<!iPendan�������!KAR�EL:*���	��KC�.�@��V�ISION SE!T���u���!�ϣ� �������	��P�'��9߆�]�o޽�CTR/L L��؃��
��FFF�9E3��u���D�EFAULT���FANUC W�eb Server��
��e�w���j��|�������WR�_CONFIG �MY�X�����IDL_CP�U_PC���B��x�6��BH�M�IN'��;�GNR_IO�K���"���NPT_SIM_�DOl�v�TPM�ODNTOLl� >��_PRTY��6���OLNK 1N�ذ�� 2D�Vh��MASTE�k�s�w�OñO_gCFG��	UO��|��CYCLE����_ASG 19O��ձ
 j+ =Oas��������//r�N�UMJ� �J�� I�PCH�x��RTRY_CN�n� ���SCRN_UP)DJ����$� �� ƣP�A��/����$J23_DS/P_EN~��p�~� OBPROC�#ܰ��	JOG�1Q�� @��d8��?� +S? /?>)3POSRE?y��KANJI_� K�l��3��#R����x�5�?�5CL_LF��;"^/�0EYLOGWGIN� q��K1�$��$LANG?UAGE X�6��� vA�LG��"S�߀�����xR��i��@<𬄐�'0u8������MC:\RSCH�\00\��S@N_DISP T��t�w�K�I��LOC��-�DzU�=#��J�8@BOOK U	L0��d���d�d��PXY�_�_�_�_��_ nmh%i��	kU�Yr�UhozoLR�G_BUFF 1-V��|o2s��o �R���oq��o�o# ,YPb���� ������(�U���D/0DCS X>u] =���"lao�����ˏݏ�3n�I�O 1Y	 �/,����,�<�N�`� t���������̟ޟ� ��&�8�L�\�n���@������ȯܯ�Ee�_TM  [d� (�:�L�^�p������� ��ʿܿ� ��$�6� H�Z�l�~ϐϢύd��SEV� ]�TYP�$���)��m�1RSK�!O�c�"�FL 1Z�� ����߯���������L	�:�TP5@���}A]NGNAM�$��E��k�UPS PG�I|%�1�%x�_L�OAD0G %�Z%CAL_T�C� ���MAXUALRM;'�I(��~���#� V�#a��CQ[x�8��n��"�t1060\	 �F�	�Ϣ����������� �� D'9ze ������� �R=va�� ������*// N/9/r/�/g/�/�/�/ �/�/?�/&??J?\? ??�?k?�?�?�?�?�? �?�?"O4OOXOCO|O _OqO�O�O�O�O�O_ �O0__T_7_I_�_u_ �_�_�_�_�_o�_,o���D_LDXDI�SAc���MEM�O_AP]�E ?=��
 �5i �o�o�o�o�o�o�o~��ISC 1]�� �oTd��\ no������ ���I�4�m��f� ��$���������!� �E�ƏT�f�:����� ß�����z��ܟA� ,�e�w�^������~� ����� �=���L� ^�2���������߿� r� �Կ9�$�]�o�(t�_MSTR ^��͂�SCD 1_xm�W���S������ �=�(�:�s�^ߗ߂� �ߦ�������� �9� $�]�H��l���� ��������#��G�2� W�}�h����������� ����
C.gR �v�����	 �-Q<u`r ������// '/M/8/q/\/�/�/�/��/�/s�MKCFG� `���/��L_TARM_2a��w2 �#�\`Y>G`METPU�T`�"����NDSP_CMNTs5p06�5�� b�΂�>�"1�?�4�5P�OSCF�7�>P�RPM�?�8PST�OL 1c2}4@p<#�
aA�!aE qOG]OO�O�O�O�O �O_�O�OA_#_5_w_ Y_k_�_�_�_�_�Q�1�SING_CHK�  +O$MODAQ73d
?�7:e�DEV 	��	�MC:MlHSI�ZEs0���eTA�SK %��%$�12345678�9 �o�egTRI�G 1e�� lf��%��?   0A$�ÜfYP�a,u���cEM_IN�F 1f>7� `)AT?&FV0E0N�}�)�qE0V1&�A3&B1&D2�&S0&C1S0}=�})ATZ�� �H�E��q9m��xAu���X�������� ������ v�)���я��П���� ���*��N����� 7�I�[�̯ן���9� &���\����g��� ��i�ڿ������ï4� �XϏ�iώ�A���m� ������߿�ѿB��� �ϊߜ�O������� �ߩ����>�%�b�t� 'ߘ�K�]�o߁���� �(�_�L���p�+����������.ONIT�OR�0G ?ak �  	EXESC1�#23E45�`789�#��x xx*x6x BxNxZxfxTrx22�2�U2�2�2�2�U2�2�2�3�3�3aR_G�RP_SV 1g��y�a(�Q>�9��?�h����?��<��@Ͽ,ѮHm�a_D�i�n�!PL_NA_ME !�5
 ��!Defau�lt Perso�nality (�from FD)� �$RR2� 1�h)deX)dh9�
!�1X d�/d/ v/�/�/�/�/�/�/�/ ??*?<?N?`?r?�? �?�?�?�?�82S/�? O O2ODOVOhOzO�O�Ob<�?�O�O�O�O _"_4_F_X_j_|_�_:LhR� 1m)9`{\b0 �_p�b�Q @D� M �Q?��S�Q?`��QaAI�Ez�  a@og;�	�l�R	 0D`4b@4c.a�P�Jd��Jd�Ki�K��J���J���J�4�J~��jEa�o-a�@���o�l[`@�z��b�f�@�S���a�Q�o�c�=��N��
������T;f�
���m[`�*  ��p  �$p>� p�$p��o?���?����������o�B ntr�Q�skse�}�l��p�  |�pu`j  #p���vks�� 	'� � ��I� �  ����}:�È~6�È=���N��b@^�d��n�Q����{�R�x���nN<. ��  '���a��`@a�@�t��@p@p�n[`C�pC0�f0�+pB�/pC3}�P��@%�Ea  �oo$|m_����gA%���. ���z�`�P���QDe���˟���(��m�� ��t O� r�u �4 ��R�c��s� :�u�a�P�` �?�ffd�!�����7� ��گ쬛af��>搠���iP�P;�e�S�_�c����>LX��s�b<	��I<g�<#��
<2��<D��<��
vo��¯��S��S.���?f7ff?u�?&찗d�@T���?��`?Uȩ?X����Z���T:z�T B��Wa�з*dů�ρ� �ϥ��������&�8�0#�\�h�+�F. K� ��G߼�3���Wɯ�����G�@ G�� ��X�C�|�g�y�� ��������jZ���� ��Q����ߙ����� 3�������/A���t_�����������d���@+Fp�IP��t��%���[`B��0����<ze�xcb!@I�
��M`B@��@�`�9@y��?��h� �@��3�[N��N��N�E��<��/:/L �>���ڟ�A�p�C�F@�S�b/�DpX������@�t��%�h���`/qG���GknF&��FצpE,8{��/ F�ZG����F�nE�DE,ڏ�/�� ���G���F7��F��ED��.��C?.?g? R?d?�?�?�?�?�?�? 	O�?O?O*OcONO�O rO�O�O�O�O�O_�O )__M_8_q_\_�_�_ �_�_�_�_�_o�_7o "o4omoXo�o|o�o�o �o�o�o�o3W B{f����� ����A�,�Q�w� b����������Ώ� ��=�(�a�L���p������(r!3�ji̹�r���ꕢ�3�㱐ڟ�y�4 �����y��P�82�D�&�jb^�p��1w����� ����ʯ���ܯ� �Js�P^�PD�c�`� m���y�\������Ӱ�¿Կ�����.� G����}ϳϡ��� 홍�U�_�J���$�y.�@�v�d�z߈ߚ� x�4�������� ��D�.�2� �$[�G�[�^�B���B��CH� ^���� u����������p�h�M�_�q�������*���^�^�Y�rm�2��
 �� ��#5GYk} ������h*��� ��>�x}���$MSKCFM�AP  ��� ����m��N"ONREL  6�9_�"EXCFENBkq
7]�FNC��}JOGOVLI�Mkduyd"K�EYk�"R�UN��"S?FSPDTYU��<v_SIGNk}�T1MOT�z�"_CE_GRP� 1n��9\ ���/���/�/4��/? �/2?�/'?h??�?C? �?�?y?�?�?�?O�? @ORO	OvO-OoO�OcO �O�O�O_�O*_<_#_�`_-�"TCOM_�CFG 1o/����_�_�_
|Q_A�RC_�6��U?AP_CPL�_��NOCHECK {?/ 5� ;h9oKo]ooo�o�o�o �o�o�o�o�o#5�GTNO_WAI�T_LF'5y"NT��Qp/���q_7ERR�!2q/_�� R_���"��:�L�dT_M�O�sr�}, ��^P_��_�PARAuM�rs/���`���MW��� =e��345678901.�@�R�)�q���_� ����˟����ݛLW��3�E�؏i�cU�M_RSPACE�,�������$OD�RDSP�SI&�O�FFSET_CAsRToݨDIS��ݢPEN_FIL�E�I!�Q�v�POPTION_IO����PWORK 5t�'� T�|�C�������䖱Z���	 �m���A�����i�_DSBL  ��v���ޡRIENTTOj���C���8=#��?�UT_SIM�_DJ�6	��V~àLCT u�}������Q��W�_PEsXE���RAT����� ���UP Sve�������ϰ���*�8��$��2��#h)deX)d�h�O�X d Y�ߑߣߵ������� ���!�3�E�W�i�{�����������2 n��)�;�M�_�q�����������<����� +=Oas����X��� O��1�m(���(��.�g��"0 ��дu�  @D��  �?��?�р��D4  E�zZ3;�	l~	 0Ӏ�S@SM� �i��i �H)!H,��H8�H�m�G�	{G�c8��6�MV��L� �C�)���)�����Ճ�*  �p  � => �  ��/�$"�,��B,�Bt�r�«����'��/���/�"��# �,0 ��� �  � �޽pj   ���&X�?MU	'� �� 12I� �  ���-�=���U?g;/�@}?�0~.ѱ�?;bѲ���H[N �?�A'M�D�> C)�f)�" B& �"O�4B+�:�Q�@�D1�oo$~����JW�AD0�J@�A: �1�E&?�O�O�#__G_2]�� ��t O� �ru �4 ���R�U��� �:�%Ёр� �?�ff��@[�_��_V_{�o~��18р"o0j>�P�Q6YPрZo�WrAdS�%��>Lw0�#�<�	�I<g�<�5�<2��<D��<�׍�l�_��ѳMb�@?f7ff?�0?&p:T�@T�q?��`?Uȩ?X�-q�iyBq5Y a��gI�_�� ����!��E�W� B�{���d�����ՏL�npΏ/�ʈG�@ G��U�ȏy�d� ������ӟ������ �yB=� ��?p���/ 򏸯�߯R���'� 9��oN�`�����~���(��ۿƿ�B�ĮD��e�ֿ;�ҿ_�J�?��h�oϨϓϸ�%�D4��b!�_@���� ߧ��Ŀ����%��@I�)�M`B�@��@`�9�@y��?�h�	� �@�3��[N��N�N�E��<�/Y��kЖ>��ڟ��A�p�C�F�@�S���pX������@�t��%�h�����!G��Gk�nF&�Fצ�pE,8{�� �F�ZG����F�nE�D�E,ڏ��ૐ��G��F7���F��ED�� Mf��b�M��q��� ���������(��8� ^�I���m��������� ������$H3l W�{����� �2VAS� w������/ .//R/=/v/a/�/�/ �/�/�/�/�/??<? '?`?K?p?�?�?�?�? �?�?O�?&OO#O\O�GO�OkO�O�O�O�N(�]�3�ji�O�a�y�	U�E3Ա��O<_�a4 ��%_7_�a�P�Q_c_ER�jb}_�_1w������]�Y�_@�_o�_1ol��P�b	Pcn~���o�O�o {_�o�oY�`��o�o ,/;M#�f0o �����Y�et� ~�i#�1�C�yM�_� ����������{bS�Ԏ���	�?�-�c�Mj2v���$�VG�z�}�B����B��CH�}�9�֟�����0�B���wl�~��������Ư�T�"��\��qQ��U
 ί�0�B�T� f�x���������ҿ�p��χ��� ��]{�x}��$PA�RAM_MENU� ?Յ��  DEFPULSE��	WAITTM�OUTl�RCV�� SHEL�L_WRK.$CUR_STYLj�;��OPT���ϧPTB����C��R?_DECSNw�Te '�!�3�E�n�i�{ߍ� �߱������������F�A�USE_PR_OG %P�%B�\��V�CCR��Ue�XÚ�_HOST !P�!�����ATt`���������|4���_TIME��� �T�  A�GD�EBUG��P�V�G�INP_FLMS�K]���TR����P+GA�� |�[����CH����TYPE
M�Y�A�;�Qz u������
 )RM_q� ������/*/ %/7/I/r/m//�/�/�/�/�/?��WOR�D ?	��	�RS��CPNS2�E��>2JO���B�TE���TRA�CECTL�PՅ�Z� a` a`{`�>q6_DT QxՅ�0v�0D������0���2��Sc�5{a�0��B���7�0�2 �0B�0B�0��2蠪�2�4�4	�4��4�4�4�4��4 ��2�4�4��4�4�4�4��4�4�4��2��4�4���2!�4"��4#�4���2&�4'��O&O8OJO\OnO �O�O�O�O�O�O�O�OR�4%X�1(�4)�4U*�4+�4,�4-�4.�4/�40 _2_D_ V_h_z_�_�_�_�_�_ �_�_
oo.o@oRodoTvb�11�42�44�4U5�46�47�49�4U:�4;�4<�4=�4�>�4?�4@�4�9 �o�o�o�o�o�o�o &8J\n�� �������"� 4��1�= �2�D�V�h� z�������¯ԯ��� 
��.�@�R�d�v��� ������п����� *�<�N�`�rτϖϨ� ����������&�8� J�\�n߀ߒߤ߶��� �������"�4�F�X� j�|���������� ����0�B�T�f�x� �������������� ,>�bt�� �����( :L^p���� ��� //$/6/H/ Z/l/~/�/�/�/�/�/ �/�/? ?2?D?V?h? z?�?�?�?�?�?�?�? 
OO.O@OROdOvO�O �O�O�O�O�O�O__ *_<_N_`_r_�_�_�_ �_�_�_�_oo&o8o Jo\ono�oV�o�o�o �o�o�o"4FX j|������ ���0�B�T�f�x� ��������ҏ���� �,�>�P�b�t����� ����Ο�����(� :�L�^�p��������� ʯܯ� ��$�6�H� Z�l�~�������ƿؿ ���� �2�D�V�h��zόϞϰ������$�PGTRACEL�EN  ��  ��������_UP y/�����������_CFG7 z�����e��<��� <��Z�l�<�$�DEFS_PD {/��a������IN'�T_RL |/����8Lԃ�IPE_C�ONFI+�}�O��<�x�WLID(�~/��?GRP 1���������@�
=��[���A?C��C
�XC)���B��r������dL�z������?� 	 r�N�8�Ҩ�� ´�����B������������A���> �6>�7�D_������� �='�=)�� ��������	B-���Q�M��� G Dz����
� �&L7p[� �����/��6/!/Z/��
V7�.10beta1�<�� B=q��"`ff@��"�>����!=�̽͏!A>ff�!@w�ff�"�\)�"D��?�  �!1@�!� �!Ap�#W��h/??*?<?K;�w����O/�?K/ �?�?�?�?O�?O>O )ObOMO�OqO�O�O�O �O�O_�O(__L_7_ p_[_m_�_�_�_��_  o�_$oo!oZoEo~o io�o�o�o�o�o�o�o� DQy{/�#F@ {yw}�y{ջy �-������/�Z? l?~?w���t�����я ���������O�:� s�^���������ߟ� ܟ� �9�$�]�H��� l�~����_ۯ��� ��5� �2�k�V���z� ����׿¿�����1� \n�j�|϶�� �����	�4�F�X�j� c�χߙ߄߽ߨ��� �����)��&�_�J� ��n��������� ��%��I�4�m�X��� ��ί����������! E0B{f�� ����H�Z� ��Vh�ϴϊ�� ��� �2�D�V�O/� s/^/�/�/�/�/�/�/ �/? ?9?$?6?o?Z? �?~?�?�?�?�?�?O �?5O OYODO}O�O�� �O�OtO�O�O_�O1_ _U_@_R_�_v_�_�_ �_�_�_"4FxBo |����o��o�o //0/B/;�__J �n������ �%��I�4�F��j� ����Ǐ���֏�!� �E�0�i��O^���N� ß՟�������A� ,�e�P�b��������� �o o2oTo.�hozo �o�����o��Ϳ�o
 گ'�֯K�6�o�Z� ��~Ϸ��ϴ������ ��5� �Y�D�Vߏ�z� �ߞ����������1� �Uy��:��� ������	���-��Q� <�u�`�r��������� ��T�f�x�n ��������� ���7"[Fj �������!/ /E/0/i/T/f/�/�/ �/�/�/�/?�//?A? l�e?w?&?�?�?�?�? �?�?�?OO=O(OaO LO�OpO�O�O����* �O_@RdZ_l_���$PLID_K�NOW_M  ~���A��TSV ��]�P�[? �_�_o�O&oo#o\o��B��SM_GRP� 1��Z� dI`~�oo$Cf~�d����D��TPbj�oLk�f�o "~�U�o>n2 T�~����� 7�4���p�D���R� ��ʏ����������6��
�T��*������QMR�c��mT�EGQK? GR��(�#��� [��/�A�S������� �����$����W�� +�=�O������������� ���S�Ͻ�S�T�a1 1��ڗ���P0� @����E�ϲ������ ���M�0�B�T�fߧ� �ߜ�����������7�P�,�m��2����N�A�<��z�3��������4���������5)�;�M�_���A6x���������7����������8(:�L��MAD  ����� ��PAR�NUM  ���Ko���SCH�
 ��
��S+UPD��xaq{��_CMP_�`� <P�z '�U�ER_wCHK����Z���RS���_�QG_MO� �%_�~�_RES_G����� ��v/{/�/ �/�/�/�/�/�/*?? N?A?r?e?w?J'��W,g/�?L%��?�?�? N#(��?OON#w�4O SOXON#��sO�O�ON#  �O�O�ON#d �O_<_N"V 1��Uua^�@cX��Pp�P_$@cW،P��P_@@cV��P�"THR_INR���pbA%d�VMASmS�_ Z�WMN�_��SMON_QUEUE ��e��`UȨ`�N�U�qN�V�2`END4a6/NiEXE]oNeW�BE\`>o/cOPT�IO;g?+2`PROGRAM %j�%1`O_�0bTA�SK_I��nOCFG �o�^9pDATAɓ�B{@ev2w��� ���z��+�=�O���s���������nzIWNFOɓ��}�!d r��!�3�E�W�i�{� ������ß՟���� �/�A�S�e�w�҇ބ���| �98q�DIT �Bׯj~WERFL~hwS~��RGADJ �^ƪA�  ,�?E��8��Q�IORIT�Y�W���MPD�SP�a�j�U�W�vT�OG��_TGp���Rj��TOE�P�1�ƫ (!�AF�PE5 ����!tcp��%��!ud�?�!�icm<�Q_��XYm_<q�Ƭ�Oq)� *������Op������������ <�#�5�r�Yߖ�}ߺ�@�߳������&�*�OPORT�a�Op�A%�_CAR�TREP~`ƭaQS�KSTA�X!*SS�AV`�ƪ	2500H809u�PT毙䕣�ƫ�����`X#�$�6�^m�URGEU`B��6A)WFP�DO�V�2��W�q�?Q�WR�UP_DELAY� �Ưe�R_HOT�hwR%z�����R_NORMAL��n��6SEMI�:y�QSKI�P���X%�x 	������� �X%-;%[m E������ �!//E/W/i///y/ �/�/�/�/�/�/?�/ ?A?S?e?+?�?w?�? �?�?�?�?O�?+O=O�OO1U�$RBTI�F��NaRCVTM쒻���m@DCRڕ���AB�
�B}�>A���@�_ݧ��{���$������V���HU����o��6���_ <	��I<g�<#��
<2��<D��<��
+__{_ �_)`���_�_�_�_�_  oo$o6oHoZolo~o i_�o�o�o�o�o�o�o  DV�_z�� �����
��.� @�R�=v�a������� ����׏�*�mN� `�r���������̟ޟ �����8�J�5�n� Y���}���ȯ����� A�"�4�F�X�j�|��� ����Ŀֿ�ӯ��� 0�B�-�f�Qϊ�m�� ���������,�>� P�b�t߆ߘߪ߼ߧ� �������(�:�%�^� A����ϸ�������  ��$�6�H�Z�l�~� ��{������������  2Vh��� �����
. @R=O�s�� ���/�*/</ `/r/�/�/�/�/�/�/��/??&?28�AGN_ATC 1��K� AT&�FV0E02;�ATDP/6/9�/2/9p8AT�A2>,AT�%G1%B960�k9+++�?,�1H�?,�AIO_TYPE  E�C/4?REFP�OS1 1� KO x�O[H/ O/�O�MNO`O�O�O �O_�OC_�Og__d_��_+K2 1� K LON_�_o�_*o�_5A3 1��_�_�_ o�o�o�o@oS4 1�Woio{o�o3W>�oS5 1��o�o�J���jS6 1�����]��H����S7 1� �(�:�t��ݏ���S8 1�����Ϗ�	���r���)�SMA�SK 1� O  q
���ɗXNO�?��1.�8�1AMO�TE  �.DN�_?CFG �U����5�0BPL_RAN�GQ�K!Y�POWE/R �Q5 a��SM_DRYPR/G %�%R����ȥTART �����UME_PR�Oׯ�d�.D_EX�EC_ENB  y�5]�GSPD=�p���Y3��TDB��洺RMÿ��MT_�ѐT��S�D0OB�OT_NAME ��S�;9OB�_ORD_NUM� ?��A/H80�0I$�_	��s	�\������ ��en��	@�}�D|���D0PC_TIME�OUT�� xD0S�232n�1�Q;� LTEAC�H PENDAN��j�5��=Q�x0�Mainten�ance Con�sK"-��"+�t4�KCL/C�}��6��|� No Use�=[߹�F���NPO�ќ�5��_���CH�_L@��U���	�J��MAVAI�L`���+��]�I�S�PACE1 2�=L ���وp��扢J@����8�?��� �� �V�w�N��������� ������4�&G
 l�}d	Q5U1����� ����`4&G
@l}d�#��2��������2 A/b/%/w/�//�/�3����	/�/-/ O/^??B?�?�?�?�?�4�/�/??&?�? J?l?{O�O_O�O�O�O�O�5�?OO1OCO �OgO�O�_�_|_�_�_�_o�6_*_<_N_ `_o�_�_�o�o�o�o�o!�75oGoYo ko}o+�o�o��� �)��>��8Rd v��H������ӏ%�F�-�[��G ;�� R�;�
�� ����ԟ ���
��.�@�����c���p���8�¯=�d ؠ��ϟ���!�3�E� W�i�_�q������x� �կ��'�9�K�]� oρ�w��ϛ���Ͽѿ ����5�G�Y�k�}� �ߡߗ��߻������w `S� @���8堯F�"�*ل�� ���߇����� �,����V�h�2�<� N������������� .L4v�R\ n�����
f�7��_MODE  y��MS ���&����Ïb���*	�&/�$CW�ORK_AD]��5��!R  ��t +/^ _I�NTVAL]����hR_OPTIO�N�& h�$�SCAN_TIM�\.�h�!R ��(�30(�L�8������! ��3��1�/@>�.?���S22��411d�8�1�1"3��@���?�?�?h���IP���@���JO\OnOE@D���O�O�O�O �O�O__(_:_L_O���4X_�_�_�8�1��;��o�� 1��pc]�?t��Di�1>��  � lS2�� 15 17oIo[omoo �o�o�o�o�o�o�o !3EWi{�� ��wc���	�� -�?�Q�c�u������� ��Ϗ����)�;� M�_���`[����ğ ֟�����0�B�T� f�x���������ү������$�7�  0 ��� om�������� ǿٿ����!�3�E� W�i�{ύϟϱ����� ��v���/�A�S�e� w߉ߛ߭߿������� ��+�=�O�a�s�� ����ߖ����� �� $�6�H�Z�l�~����� ���������� 20DVP�\�  �A� ������ %7I[m��������/ �/C(/N/`/r/�/ �/�/�/�/�/�/?Fa;/?B?F�x1� ;?w=	12345678{_��l�@�P�?�?�?�?�?O9/2ODOVOhOzO�O �O�O�O�O�O-/
__ ._@_R_d_v_�_�_�_ �_�_�O�_oo*o<o No`oro�o�o�o�o�_ �o�o&8J\ n���o���� ��"�4�F�X�j�|� �����ď֏���� �0�B�T�f������� ����ҟ�����,� >�m�b�t����������ί����(��6 yI�[�@�`����������Cz  Bp�*   ���2�54F��$SCR_�GRP 1�(��e@(�l���0@ >`1 [1s�	  )�3�C�<�t�vrY��8P�}�kϤ���-�95C����-u���ȡ���LR� Mate 20o0iC �190�1�Շ0LR2C ��3�=OÆ�D�
f؜1u�2�U7��`1���v��@�u���	�t���������$�^0�2���_2T�g� �ϊ��o�F�D�f?��s�����￶ht ,oZ�k`r�B�˰!�P�N�g�N�Aܰv�G  @DЎ�N�@�����  ?� ��J�H�˰��y�N�F@ F�`������ A,Qwb��� n�N�������B��_J� n�����/� %//I/��E+:3��6?|?�5��
�/�/�#��=@=��"�/p�l�� 3B�07�5�90@7���EL_�DEFAULT � I����� ^1MIPO�WERFL  �V�v5]2�0WFDO�k6 v5 �ERV�ENT 1����O�t3C�L!DUM_EIP?��8�j!AF_�INEj0O�$!�FT�?=NOaO!�Q�O �PO�O!�RPC_MAI�N�O�H��O�O�CV�IS�O�I��OE_!7TP8PPU<_�9�d4_�_!
PMON_PROXY�_��6e�_�_XR�_�=f��_)o!RDM_'SRV*o�9gouoG!RR8�o�4hdo��o!
�@M�_�<i��o!RLSY3NC4y8�oY�!ROS�?�|�4H�tO�8c�� ���;��_�&��� J���n������ȏ ڏ7�I��m�4���X�����7ICE_KL� ?%�; (%�SVCPRG1@�����!��3*�D/��4R�W��5z�D��6�����7ʯ ϯ�C��5�9��oG����o�� ����D����l�� 񑔯�񑼯7��� _������4���� ]�����������'� �տO����w��%� ���M����u���� ������?�A��Ͽ� ђ�؟ꐊ���ɱ�� ������?�*�c�N� �������������� ��);_J�n ������% I4mX�|� ����/�3// W/i/T/�/x/�/�/�/ �/�/�/?/??S?Ś_DEV �9��MC:[8�wim4OUT_R�f1~6i8REC �1���f0�0 �f0 	 f0.�2  
f0�4�1 ���3OMK�1�4�=A%O^OAA��
 ��Z�6 s ;B�3AAqE=�=A���2TWG�1f0)f0{f0�U�Of2B0�����/Q0�O_�5T��@��@r�H�;@_�  x�0}@�U@��O f0��f4�1af0�V_�2X�0��@�f0?�@�X~_�__��2\�0���0��0�@��-��_ f0�f0�1�=f0[f0�o�2T�0��@�f0*�@uX*oco�_�ÆLH�0��0��R � G �RobmU�f0Ezf0�o�2�Q��@�f06�@z�ovo�~K�L=A�1(f0t"f0�f0�_c�f4e�Z=�ZZ f0k0U��0Cf0f0q��"~N�LiI�1�2�f2Pf0>jI��zDf0f0o.�g����φL"f0i�0b*f0��0��0V�bU�f0f0/f0|~S 0��E0��@�f0$�@Y�^�p����ՆL*�A�0=�Qp�ɀ��b�ʈ�Rf0_^�f2C0��@���A0����&���2\�AM��Up��A��p�<~��O���Ӧ�$2�k�ҟ��2\&f0}��0J�0Wf0�Z��b�f0�f0R~�[���F��@ݒq0"ޯ�*� a@��Z�H�~�l� ������ؿ������ 2� �V�D�zό�nϰ� ������������.�� >�d�R߈�v߬ߚ��� �������*��:�`� N��f�x������� ���&�8��\�J�l� n������������� ��4"XFh�p ������0 B$fT�x��x���5V 1��<���`��A!O  _ -�P��}�a?_TYPE�?�k2HELL_CFOG �z:f2/� HL�/<7RS ա�/�/�/"??F?1? j?U?�?y?�?�?�?�?��?O�?0OBOQK�
�p�!%QOO�O%���x�q�qQ��M�q�p�$�gBQ�d�O�O�&�HK 1��+ �OE_@_R_d_�_�_ �_�_�_�_�_�_oo *o<oeo`oro�oa&�#?OMM ��/�o��"FTOV_EN�M�t"!}*OW_R�EG_UI�o�"IMWAIT�b���G.${OUTv$&ywTIMu��`�VAL5's_UN�IT�c�v})MON�_ALIAS ?�e�i ( he !� ��$�6�%�� c�u�����D���Ϗ� ����)�;�M�_�q� �������˟ݟ��� �%�7��H�m���� ��N�ǯٯ������ 3�E�W�i�{�&����� ÿտ習���/�A� �e�wωϛϭ�X��� ��������=�O�a� s߅�0ߩ߻����ߊ� ���'�9�K���o�� ����b�������� #���G�Y�k�}���:� ����������1 CU y���� l��	-�Q cu�2���� ��/)/;/M/_/
/ �/�/�/�/�/v/�/? ?%?7?�/[?m??�? <?�?�?�?�?�?�?!O 3OEOWOiOO�O�O�O �O�O�O�O__/_�O @_e_w_�_�_F_�_�_ �_�_o�_+o=oOoao soo�o�o�o�o�o�o '9�o]o� ��P�������s�$SMON_�DEFPRO ����:�� *SY�STEM*  ��l�*�RECA�LL ?}:� �( �}7cop�y virt:\�output\c�alprz.pc� md: ove�r =>1014�49728:95?1961  ����a3�Џ⏻p}8z���tcp������D��V��:����_dv?_xy.ls���5�Ɵ؟�Fz�����tp~������A�S�&e�}9z���z����P4�ůׯ�D��z� �����A�S�e�����������3�Ŀֿi��tpdisc 0�=>laptop�-3jv248m�s:20980 �������O�a�t�t�pconn 0 ���'�9�����o�
�xyzrate  ���ϗϩϻ�L�^�q��!���13960 �.�f�����v�y������372244�48:87818C5 ��C�U�h�A�� �����-�<�����2r�5���_1�"�@��A�S�e���
�2� #�5���������ޠ� ��CUh�z�0 �����
���� DVi�{��!�0� ��������&��I/[/n�6���/ �1/�/�/g/�\test��"/�/E?W?j� ��5��8?7?�?�? m/�?����?DOVOi�?z:	��GO�<O�O �Or��O&�OE_W_j�E�����"��_�_ �_w����_,�_DoVo�]C���_��O�o�o �o�/�o��oOa t��3��i {����B�T���o ��/��ҏ�w�o@��!���O�a���;z��frs:orde�rfil.dat��dtmpback�\��6�ǟٟlZ2>zTb:*.*����@�Э��P�b��2xz�:\�����1�¯ԯg�7z�a������ ��C�U�h�z����0� ��ӿ��������?��Q�c�  �$SN�PX_ASG 1߶������� P 0 �'%R[1�]@1.?_��?�pS%���Ͽ� ����� 6��@�l�Oߐ�s߅� �ߩ������� ��� V�9�`��o���� ���������@�#�5� v�Y������������� ��<`CU �y������ &	0\?�cu �����/�/ F/)/P/|/_/�/�/�/ �/�/�/?�/0??%? f?I?p?�??�?�?�? �?�? O,OOPO3OEO �OiO�O�O�O�O�O�O _�O _L_/_p_S_e_ �_�_�_�_�_ o�_�_ 6oo@oloOo�oso�o �o�o�o�o�o  V9`�o��� �����@�#�5� v�Y�������Џ��ŏ ���<��`�C�U� ��y���̟���ӟ� &�	�0�\�?���c�u� �������ϯ����F�)�P�|�_�x�PA�RAM ���}�� �	����P��p�OF�T_KB_CFG�  ����״PI�N_SIM  ��̶�/�A�ϰx��RVQSTP_DSB�̲}Ϻ����SR �	�� �& CAL_T�Cŵ�Ͻ�ԶT�OP_ON_ER/R  ������PTN 	���A��RI�NG_PRM�� ���VDT_GR�P 1�����  	з��b�t߆ߘ� �߼��������+�(� :�L�^�p����� ������ ��$�6�H� Z�l�~����������� ���� 2DV} z������� 
C@Rdv� �����	/// */</N/`/r/�/�/�/ �/�/�/�/??&?8? J?\?n?�?�?�?�?�? �?�?�?O"O4O[OXO jO|O�O�O�O�O�O�O �O!__0_B_T_f_x_ �_�_�_�_�_�_�_o o,o>oPoboto�o�o �o�o�o�o�o( :Lsp���� ��� ��9�6�׳�VPRG_COUNT�����d�'ENB/�_�M������_UPD 1�>	�8  
M��� ����-�(�:�L�u� p���������ʟܟ�  ��$�M�H�Z�l��� ������ݯد���%�  �2�D�m�h�z����� ��¿Կ����
��E� @�R�dύψϚϬ��� ��������*�<�e� `�r߄߭ߨߺ��������\�YSDEBU)Gn�Ӏ� �d��"�SP_PASSn��B?4�LOG [�΅�� �9��
�  ��� �?
MC:\`��a�_MPCf�΅��$��ҁ��� ҁ��SAV �i�؆�� ���SV��TEM_TIM�E 1�΋ (�J��F�}��%��T1SVGUNSɀ�o�'�����AS�K_OPTION�n�΅������BC?CFG �΋O�c H�2!`; A�I�r]o��� ����8J5 nY�}���� �/�4//X/C/|/g/�/�/ ��,�/�/  ??�/�/H?3?l?W? �?��?��0�?�?�? O�?&OOJO8OZO\O nO�O�O�O�O�O�O_ �O _F_4_j_X_�_|_ �_�_�_�_�_o�X�   o2oPoboto�_�o�o �o�o�o�o�o: (^L�p��� �� ��$��H�6� X�~�l�����Ə��� ؏�����D�2�h�o ������ԟR���� �.��R�d�v�D��� �������Я���� <�*�`�N���r����� ��޿̿��&��J� 8�Z�\�nϤϒ���~� �����"�4߲�X�F� hߎ�|߲����ߤ��� ����B�0�R�T�f� ������������� �>�,�b�P���t��� ����������(�� @Rp���� ���$6Z H~l����� �� //D/2/h/V/ x/�/�/�/�/�/�/
? �/??.?d?R?�?> �?�?�?�?�?r?OO (ONO<OrO�O�OdO�O �O�O�O_�O__&_ \_J_�_n_�_�_�_�_ �_�_�_"ooFo4ojo Xozo|o�o�o�o�o�?  0BT�oxf �������� �>�,�b�P�r�t��� ������Ώ��(�� 8�^�L���p�����ʟ ��ڟܟ�$��H��o `�r�������2�دƯ�����2��P��$�TBCSG_GR�P 2����  �P� 
 ?�  {� ��w�����տ��ѿϠ��/�A�T�[��b�_d0 �p�?P��	 HBHA�L��͌�@�B   C����϶ˀ��ϟ�D�����A���x���A���T$�9��6ff���f�@P�C�ώ�@1�f߬��C��ߐ� �ߴޥ���%��%�D� W�"�4���j�|�������?Y������	V3.00~s�	lr2c��	*2�*�O�A� �.�ѳ33P�d���� x�J�y�  �������T�JCFG� ��l� �o�����������=K
 %�Kq\���� ����7"[ Fj����� ��!//E/0/i/T/ f/�/�/�/�/�/�/s� ��??(?�/[?F?k? �?|?�?�?�?�?�?O !O3O�?WOBO{OfO�O �OP�<��O��O�O�O 0__T_B_x_f_�_�_ �_�_�_�_�_oo>o ,oNoPobo�o�o�o�o �o�o�o:(^ L������h�  ��$��H�6�l�Z� |�����Ə��֏؏�  ��D�V�h�z�4��� ����ҟԟ��
� @�.�d�R���v����� ���Я���*��:� <�N���r�����̿�� �޿ �&��>�P�b� ϒπϢϤ϶����� ���4�F�X�j�(ߎ� |߲ߠ���������� �B�0�f�T��x�� ����������,�� P�>�t�b��������� ������&(: p^����t�� ���6$ZH~ l������� /2/ /V/D/z/�/�/ �/j/�/�/�/�/?.? ?R?@?v?d?�?�?�? �?�?�?�?OO<O*O `ONOpO�O�O�O�O�O �O_�O__&_\_� t_�_�_B_�_�_�_�_ �_"ooFo4ojo|o�o �o^o�o�o�o�o�o 0B�oxf�� �������>� ,�b�P���t������� ��Ώ��(��L�:� \���p�����ʟ���  ��_�*��_�l�Z� ��~�����į�د�  �2���h�V���z� ��¿Կ濠�
���� �.�d�Rψ�vϬϚ� �Ͼ������*��N� <�r�`߂߄ߖ��ߺ� ������8�&�H�n� \���>�����x�� ����4�"�X�F�|�j� ��������������
 Tfx�D� ����� P>tb���� ���//:/(/^/ L/n/p/�/�/�/�/�/  ?�/$?6?��N?`?r? ?�?�?�?�?�?�?�?  OODOVOhOzO8O�O��O�O�O�O�N  PS V$_R��$TBJOP_�GRP 2��E��  �?�W<RCS�J\=��@0WP�Ry@T�P � ��T��T �Q[R	� �BL  �UCр D*W[Q�_��_?fffe:�lB �P�ff�@`�33D  $a�U3o>g�_�_�po�l�P�e9<�b>bY��?٪``�$o�oUA��gD�`$�co�Quz�9�P�Aa�P@>a���C�Z`Ep<�o]A6ffpu`asD/�U�h�͔r ��~�a�RieAq�`�q���@9q�|�d&p`%���c333D��\P8���?�`?1L�pAp[QB�b�k��}� ��z�� >�sffԁL���T� f��fo ��Nw@�*� 8�f���r�,���П�� ȟ��'����F�`�J��X�����SC�V�ء��	V3.0}0�Slr2c�T�*��TQ��� E���E��A E��E���3E�iNE��!hE�فE����E�I�E���E���E��rF�F��FM(F��5FBF�aOF�\F"�f,�z  E��@ E�� E��� E�  E������ E������ EȆ�Ԏ������ F   �F� F$ �Fj` F�@ �F�P F�` �9�IR9�o���L�_ ��V��LQ�8TESTPARS��XUP9SHRk�AB_LE 1�J[4�SV�+� �0�VǅV�V�WQV�	�V�
V�Vȥ�Q�V�V�V�뱅�RDI��TQ�϶���������f�On߀ۊ� �߮����ކ�Sl�RS 0ړ��������� ���#�5�G�Y�k�}� ������������/]k� o��*	�%�7�I��π��+�=�O؆�N�UM  �E*TQ�PP �����_CFG �����Q@<PIMEBF_TTq��RS~�;VER�<Q�;R 1�J[
' 8�RP� �@5  ��� ���//&/8/J/ \/n/�/�/�/�/�/�/ #?�/?Y?4?F?\?j?�|?{_�h@R
�<PMI_CHAN�G R �3DBGLVQ`IR;Q�0�ETHERAD �?�E;@�S ��?�?TO6V�0ROUmTe!JZ!�D��OwLSNMASK�0HRSAA255.��E��O�O8TOOL�OFS_DIq���5IORQCTRL �s[���n]8]_�_�_�_�_�_�_ �_o"o4oFo�
�_To�fo�og�PE_DE�TAIH3ZPON?_SVOFF)_�c�P_MON ��"P2�iSTRT�CHK �J^�mO�bVTCOMP�AT�h;C�d�`FP�ROG %JZ%�  AL_TCPx=�n%QPLAYr���j_INST_M��@ �|�g�tUS8e]orLCK��{QUICKME�0�)�orSCREF�}3Jtps��@or�a�f��2w�_{����ZyISR_GR�P 1�JY ؛ 6���@��;�)�_�M��8 ����Y�������͕ �����/��S�A�w� e�������ѯ��������=�+�M�s�	�12345678h����f�X`�1�Ћ�
 �}ipn�l/۰gen.htm�����0�B��X�Panel� setupF�}�<�ϘϪϼ����� u�k��*�<�N�`� r��ϖ�ߺ������� ��ߝ�J�\�n�� ����I�?������ "�4�F���j������ ��������_�q�0 BTfx��� ����>� bt����3�~�UALRM�pG {?J[
  � */!/R/E/v/i/�/ �/�/�/�/�/�/??�<?�SEV  ��n6�ECF�G ��m�6��A��1   Bȩt
 =?�s3E�?�?�? OO+O=OOOaOsO�Oh�Gz1ʂ��k S(Ο�OH7Isv?}{�`(%0?"_p_I_4_ m_X_�_|_�_�_�_�_��_o�_3o�L� ��M�OAoI_E�HI�ST 1��i  �( k`���%/SOFTPA�RT/GENLI�NK?curre�nt=editpage,,1 �q��`�o�o'z�(��o�emenu�b955�`�ou��(�:L148,2 _XYd�� ��,��}53�aZ�� ����2�D��0n�����"�4�À'ǏM~3	4�`�`4�����r��,K��nCAL�o���*�<�G�Y��`71�`MV��������í�)a�a)o��� %�7�I���ޯs����� ����Ϳ\����'� 9�K�ڿoρϓϥϷ� ��X�j����#�5�G� Y���}ߏߡ߳����� f�����1�C�U��� �ߋ���������Я 	��-�?�Q�c�u�x� �������������� );M_q �� �����%7 I[m��� ����!/3/E/W/ i/{/�//�/�/�/�/ �/?��/?A?S?e?w? �?�?�/�?�?�?�?O O�?=OOOaOsO�O�O &O�O�O�O�O__'_ �OK_]_o_�_�_�_4_ �_�_�_�_o#o�_Go Yoko}o�o�o�oBo�o �o�o1?�og y�����o�� 	��-�?��c�u��� ������L�^���� )�;�M�܏q������� ��˟Z����%�7� I�؟��������ǯ ٯh����!�3�E�W��Bz�$UI_PA�NEDATA 1��������  	�}�/frh/cg�tp/wided?ev.stmc����ҿ����)pri��.�Ip}2�V�h�0zόϞϰ� )���� �������0��T�;� xߊ�q߮ߕ���������Bv�� �(� # Q� @�E�W�i�{����� ��6�������/�A� ��e�w�^��������� ������+O6 s�l�� ��� ������1C �g������ �L	///?/&/c/ u/\/�/�/�/�/�/�/ �/?�/;?M?���? �?�?�?�?�?0?Ot %O7OIO[OmOO�O�? �O�O�O�O�O_�O3_ _W_i_P_�_t_�_�_ �_�_Z?l?o/oAoSo eowo�_�o�o O�o�o �o+�oO6s �l������ �'�9� �]�D����_ o�oɏۏ����#� v�G��ok�}������� ş,�������C� U�<�y�`�������ӯ ����ޯ�-�����c� u�����������T� ��)�;�M�_�q�ؿ ��|ϹϠ�������� ��7�I�0�m�Tߑߣ� ����:�L����!�3� E�W��{�� ϱ��� �������r�/��S� e�L���p��������� �� =$a����}�r�����)�*��V hz����� ���.//R/9/v/ �/o/�/�/�/�/�/?��������$UI_�PANELINK� 1����  �  ���}1234567890_?q?�? �?�?�?�4��]?�?�? OO1OCO�?gOyO�O �O�O�OYIY0:�M���[0-/SOF�TPART/GE�NA1?CONFI�G=SINGLE�&PRIM=mainedit �O�I_[_m_YJ_$_M=�wintpe,1`@_�_�_�_XK  �_ $o6oHoZolooo�o �o�o�o�o�o�o
2 DVhz��� �����.�@�R� d�v��� �����Џ�����M 0,mM9P E=Por?>S�,Ico:�{� ^�������˟ݟ��� ��7��[�m�P������O���BS0ߢ��C���/�%�7�I� [�m�`C�������Ϳ ߿񿀿�'�9�K�]� o��L���э͙�Q|� ���������!ߨ�;� M�_�q߃ߕߧ�6��� ������%��I�[� m����2������� ���!�3���W�i�{� ������@������� /��Sew�� ��.���z�! E(W{^�� ����/�//A/ ���͡Ϸ�}����/�/ �/�/�/?�2?D?V? h?z?�??�?�?�?�? �?
OO�ϝϯ�dOvO �O�O�O�OE�O�O_ _*_<_N_�Or_�_�_ �_�_�_[_�_oo&o 8oJo�_no�o�o�o�o �o�oio�o"4F X�o|����� e���0�B�T�f� ���/��������� ُ���>�P�3�t��� i�����Ο��O/�s/ (��/L�^�p������� ���?ܯ� ��$�6� ůZ�l�~�������#O 5OGO�� �2�D�V� h���Ϟϰ������� u�
��.�@�R�d�v� ߚ߬߾������߃� �*�<�N�`�r��� ������������&� 8�J�\�n�������� ��������m�"4ß XjM�q��� ���BT7 x������A�� //,/>/P/C�t/�/ �/�/�/�/�/o/?? (?:?L?^?Ϳ߿�? �?�?�?�? OO�?6O HOZOlO~O�OO�O�O �O�O�O_�O2_D_V_ h_z_�_�_-_�_�_�_ �_
oo�_@oRodovo �o�o)o�o�o�o�o *�oN`r�� ���m��&� 8��\�n�Q���u��� ȏ������"���?��?�{��$UI_�POSTYPE � �5�� 	k�{��_Q�UICKMEN � ��j�����RE�STORE 1���5  ��/
�2�D�h�mc�������¯ԯw� ��
��.�@��d�v� ������W���˿ݿO� �*�<�N�`�τϖ� �Ϻ����ρ���&� 8�J���W�i�{��϶� �������ߡ�"�4�F� X�j��������� �ߋ����y�+�T�f� x�����?��������� ��,>Pbt� ����� (�L^p����I��� //��S�CREܐ?��u1sc-��u2M$3M$4M$5*M$6M$7M$8M!���USER/ 4/F"TL. O#ksW#�$4�$U5�$6�$7�$8�!���NDO_CFG� ؜�  ,� ���PDATE ��)�No�ne V��SEU�FRAME  �
��&,1RTOL_ABRT7?��N3�ENBX?I8GRP� 1�!��Cz  A��3�1��? �?�?�?�?FO"O�G:ېUx81g;MS�K  {5�Ag;N&41%a��B%��O���VISCAND�_MAXyEI��c8�@FAIL_ISMGy@f���#�8��@IMREGNU�MyG
�KRSIZlyC,���$,S?ONTMOUW0{D��%�VU�#�cװ� �P�2�FR:\�O � MC:\XS�\LOG�VB@4 !�O�_�Q�_o�
�z MCyV�_�SUD10fEX9k
�f�wV�2�ۜ��p(��=��͓o��j�o�o �o�o�o�o�o 2�DVhz��KPO�64_?S�0��3n6�uQ0LI Q�z��x�qV� �|f@��w�� =	�xS�ZV�~����wW�AI��DSTAT' ܛ;�@�_ď�֏�$����EP12�DWP  ��P G/����q�AP�-��B_JMPER�R 1ݜ�
  �� 2345678901�������ʟ ��ϟ��$��H�;��l�_�q����LT@ML�OW���P�@�P_T�I_X�('�@MPHASE  5�3��CSHIF�TUB1~k
 <���Ob��A�g��� w���ֿ�������� �T�+�=ϊ�a�s��� �ϩ��������>�ߠ'�t�K�!��#ޛ:	�VSFT1�suV�@M�� �5���4 �0��UA� W B8���Ќ�0p�����Ҫ��e@��#ME*�{D�'���q���&%�!�M�$ߴ~k��9@�$~�T?DINENDcXdH�z�Ox@[O��aZ��Sp����yE����G����2������x����RELE��y?w�^_pVz�_AC�TIV���H��0A ��K��B#&���RD�p��
1YBO�X ��-�����2�D��190.0.� 8�3��254��2�p�&���rob�ot�ԟ   �pN g�pc� �{�v��x���$%ZABC
�3�=,{�낆 ;-!/^/E/W/i/{/�/ �/�/�/�/?�/6??H/?l?!ZAT����