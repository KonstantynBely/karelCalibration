��   ?3�A��*SYST�EM*��V7.7�0107 10�/3/2018 A   ����MN_MCR�_TABLE �  � $MA�CRO_NAME� %$PRO�G@EPT_IN�DEX  $OPEN_IDa�ASSIGN_T�YPD  qk$MON_NO}�PREV_SUB�y a $USER�_WORK���_�L� MS�*RT�N  &S�OP_T  �� $�EMG�O��RESE�T�MOT|�H�OLl��12��STAR PD�I8G9GAGBzGC�TPDS��REL�&U�s �� �EST�x��SFSP�C���C�C�NB��S)*$8�*$3%)4%)5%)6�%)7%)S�PNS�TRz�"D�  ��$$CLr   O����!������ VIRTUA�L�/�!;LDUI�MT  �������$MAOXDRI� ��5��%.1 �%� � d%�Open han�d 1����% ta?�? �"  �!��#q0Close�Q?d?�?�?�9�7Relax�?�?)OOO�9�6L82QO2O�O VO�3 �?�O�O
_�O�4O�O�Ol__�6�Fh_�_d_�_�[�3 ��
@�_o�_<o�_�_ ro!o�o�oWo�o�o�o �o�o8�o5n /�S�w��� �4���j����=� O���֏��������0� ߏT���O���K��� o��������,�۟� b����5�G���k��� 򯡯��(�ׯL���� �������g�y�� ���ӿ�Z�E�~�-� ?ϴ�c��χϙ��� � ��D����z�)ߞ߰� _ߙ��ߕ�
����@� ��=�v�%�7��[��� �����<����� r�!���E�W������� ����8��\ W�S�w��� "4�j�= O�s����0/ �T///�/�/�/�/ o/�/�/�/?�/�/? b?M?�?5?G?�?k?�? �?�?�?(O�?LO�?O �O1O�O�OgO�O�O�O _�O�OH_�OE_~_-_ ?_�_c_�_�_�_o o oDo�_ozo)o�oMo _o�o�o�o
�o�o@ �od%_�[� ���*�<��%� r�!���E�W�̏{�ɏ ���Ï8��\��� ������ȟw������� "�џ��j�U���=� O�įs�诗����0� ߯T�����9����� o��������ɿۿP� ��Mφ�5�Gϼ�k��� �ϡ��(��L���� ��1ߦ�U�gߡ����� �����H���l��-� g��c�������� 2�D���-�z�)���M� _�������
����@ ��d%���� ��*��% r]�EW�{� ���8/�\/// �/A/�/�/w/�/�/�/ "?�/�/X??U?�?=? O?�?s?�?�?�?O0O OTOOO�O9O�O]O oO�O�O�O_�O�OP_ �Ot_#_5_o_�_k_�_ �_�_o�_:oLo�_5o �o1o�oUogo�o�o�o �o�oH�ol- �������� 2���-�z�e���M� _�ԏ���������@� �d��%���I���П ������*�ٟ�`� �]���E�W�̯{�� ����&�8�#�\��� ��A���e�w������ "�ѿ�X��|�+�=� w���s��ϗϩ�����B�T��=�
Send EventU��5�SENDEV�NT��3�i�� %	}�Data<�ߘ�DATA�߿����%}�Sys�Var��SYS�VY��1�%G�et��Z�GET�����%Re�quest Me�nu����REQM'ENU!�����?� ��;ߤ�_�������� ����F��j+ �O����� 0��fxc�K ]������>/ )/b//#/�/G/�/k/ }/�/?�/(?�/�/^? ?�?�?C?}?�?y?�? �?�?$O�?!OZO	OO �O?O�OcOuO�O�O�O  _�O�OV__z_)_;_ u_�_�_�_�_�_o�_ @o�_o;o�o7o�o[o mo�o�o�oN �or!3�W�� ����8���n� ��k���S�e�ڏ���� ������F�1�j��+� ��O�ğs�������� 0�ߟ�f������K� ��ү��������,�ۯ )�b��#���G���k� }����(�׿�^� ς�1�C�}��ϵ��� �ϯ�$���H���	�C����?ߴ�c�u��$M�ACRO_MAX�:�������Ж��SOPE�NBL �����՗�r�r�A�����PDIMSK�����Y�SU�c�u�TPDSBEOX  -�q�U����n����