��  ë�A��*SYST�EM*��V7.7�077 2/6�/2013 A�Q  �����ABSPOS_G�RP_T   � $PARAM  ����ALRM_RE�COV1   �$ALMOEN5B��]ONiI �M_IF1 D� $ENABL�E k LAST�_^  d�U��K}MAX� $LDEBUG@ � 
GPCO�UPLED1 �$[PP_PRO?CES0 � ��1�FPCURE�Q1 � $�SOFT; T_I�D�TOTAL_�EQ� $,N�O/PS_SPI�_INDE��$�DX�SCREE�N_NAME {�SIGNj���&PK_F�I� 	$TH{KY�PANE7�  	$DUM�MY12� �3��4�GRG_S�TR1 � �$TIT�$I��1&�$�$T�$5&6&7&8&9'0''��%!'�%5'1?'1*I'1S'1]'2h"GSBN_CFG1 � 8 $CNV_JNT_* ��DATA_CM�NT�!$FLA�GSL*CHEC�K��AT_CE�LLSETUP � P� HOM�E_IO� %�:3MACROF2R�EPRO8�DRUeNCD�i2SMp5�H UTOBACK}U0 � �	�DEVIC#TI\h�$DFD��ST�0B 3$INTERVAL��DISP_UNI�T��0_DO�6E{RR�9FR_Fa��INGRES��!Y0Q_�3t4C�_WA�4�12HGX�_D�#	 d �$CARD_E�XIST�$FSSB_TYPi�� CHKBD_S�E�5AGN G�� $SLOT_�NUMZ�APRE�V��G �1_E�DIT1
 � Uh1G=H0S?@�f%$EPY�$OPc �0L�ETE_OKzBU�S�P_CRyA�$�4�FAZ0LACIwY1KR�@k �1�COMMENy@$DGV]QP� h���AL*OU�B? , $�1V$1AB0~ OL�U=R"2CAM_;1� x�f$A�TTR��@0AN�N�@�IMG_H�EIGHyAcWI7DTH�VTCYU��0F_ASPE�CyA$M@EX�P;$� Mf�C�FcD X $�GR� � S!1U`BfPNFLIC`~d
�UIREs3��AO}MqWITCH}cJX`N.0S_d�SG0� � 
$WARNM'@f��@� sLI? �aNST� �CORN��1FL{TR�eTRAT@0�T�`  $ACC�1"p '|�'r�ORIkP�C�kRT�q0_SF� O��CHGI1� [ Tz`u3I�PpTYVD�@*2 ��P�`� 1zB*HED�SJ* ��q2�vU3�v4�v5�v6�v�7�v8�v9�CO�$ <� so�o�h��s1�PO_MOR~. t 0�Ev�NG�8`TBA� 5c���A�����]@����ϋaP�0Ѕ*��h�`
P�@�2� �,p�J,p_Rrrqo@+�1J/r/�J�JVq@�Cj��m�g��usp�q�P_}0OF� 2 ; @� RO_����WaIT8C��NOM	_�0�1ەq3W ��cD �;����hP���mEXpG�0�� F�p%r
$T�Fx�JF�D3ԐT�O�3&@U=0�� ��H�24�T1��E�� �e��f���f��0CPDBiG;a� k@$�P�PU�3�f)�:��A�AX 1�dU�N�$AI�3BUFpuF����! |�`l��`PI��Pr�Mq�M~�䠁�}Fr�SIMQS���G��QE�����_M�C{� �$}1JqB�`S�}1DEC��౐��(�?�z� ���0CHNS_EMP�r$Gg�=Ǎ@�_��q3
p1_FP󔞡TCh�@`�b��@q0�c}�y�G�� V�A0Ԃ�!!���JR!0Ԃ?SEGFRA.pv �7aR�T_LIN�C��PVF������Y���Q���)B����( ' ���f�e�S���Q��.0��p�B��A����SI!ZC�ћ�z�T��g�������QRSINF 3��p����?�������؉���Lot��G�*�gCRC�eFCCC�` +���T�h��mh�SbA@��h�*�f��:�D�dd�c��C��PTA��`��w@�撀��EV���jF��_��F��N�&�G�� X�������1i��! ��,��hRGNP��0qF���R}�D���2}�LEWN��Hc6����C�K�(�RcDx :�L��ou2���A�6N`Co�$LGp��B�1aP��s@�dBWaA?@���~0R����dME%`��d�f_RAs3dAZCh���z�OkqFC�RH`X`F�`��}��,�ADI;� 6b � ���`�p�`5cn�aS�@1�7a�AMP����PY8CU�M��CU��iQU� $�P��C�CG1�������DBPXWO�����p$SK���2۱DBT TKRL�1 ��Q0Ti�� �P�DJ�4LAY_CAL�1R �!'PL	3&@�0EAD�Q5'�Q5'̡�d��1!�W�PR� 
�1 0�1"� �PA$�q�$�� �L�)#��/�#mp�0$�/�$Cr�!%�/�$ENEq�r�&�/�#d RE|p�"'H ��O)@"$LF3#�$�#xB� W;���FOf[ _D0m�RO(@����u��j���3RIoGGER�6PA%S|���ETURN�2nRcMR_��TU�`�?�u0EWM��Ƹ�GN�P��zBLAx��E��$$P#�CP� ��&@�Qk�C5D�mpD�A#�p4�\1i�FGO_AWAY�2MO��fQg��CS_(<�QIS ���@�c�C���A����B@�t�Cn��A"�FW��N�DNTV@��BVkQ������S˳W�sU�J�&�U�� ��SAFE��ZV_SV6bEX�CLUl�����ONLA��SY��Q�t�OTBa��HI_V|/M�PPLY_�a>��VRFY_#�qx�Bd�_ )0����_+�Ip ��TSG3� * �b݀�0 AM���a*�����0��Vi.b%fA�NNUN� rLdI%Dp�U�2~S@�`�mijarj�f�pO�GI�"+��$F�Ob�׀OT@w1� $DUMMY ���d[!�d١�& ��E, ` 8�HExs��b�SB$��SUFFI��@ ��@�a5�g6��a�MSW�E- =88�KEYI���ÃTMZ1^ӌq�1�vI�N�����. �D��HOST? !�r���t[ �t٠�tYp�pEM>���$���SBL��UL��/� �|3����T�50�!0 � $<9��ESAMP�ԕ F��������I�0�>�$SUBe�Q��� �C�:��G�SAV��r���G�C� ˇ,�PnfP$80E���YN_B�1 0&�`DIad�@O���v}$]�R_I��� �ENC2_	ST � 2
ԇ J���L�q~S�`;����!!3�M�I��1:�p�4  L�3�M���0�0K�4'a��A�VER�q��}�M�D3SP�v��PC�U����\ì�VALMUŗHE� ��M�sIP@���OPP7  �THS ���6��S�F�F􁳠d0L�0�T��SC�Q�dm:�ETo�5zrFULL_DUY��da�0��O�w�h�O�T���0NOAUkTO�!6�p$�H\���cl�
�C��%�C�������L�� 7H *�L���n�b���$�0P�˴��ֲ��[!����a��Yq��dq��7*��8��9��0����U1��1��1��1ȺU1պ1�1�1���2
�2����2��2���2Ⱥ2պ2�2��2��3
�3��3T����3��3Ⱥ3պU3�3�3��4
��)[���SE�"8 A<��~��`�;I��0���/��QFE�0�0�� 9 ,��Q?3 z@^ ?�А
��ER@#����A��� :�`$TP~�$VARI��<��UP2�P; �pq�TD��S|�1`�3���e�BAC��< T�pr��)��bP�P o�IFI@)�P ���U���P���P��0��� =t� ;'�Ԡ��P'�ST(&�� HR&�r0E�T���	%�C��	� ��_Cr�N�r��B��p��h�FORCEUP�%bn�FLUS�`H�N �E�h�RD_�CMK@E(����I�N_��&vPg�REMM�F~Q��M ��( 3
K	N0��EFF��N@IN��A��OVMl	OV=Al	TROV����DT��mDTMX ���m{@�
��? ��*[ ��CL��_ :p']@$�-	_
�;�_T��X
��@AQD� ��}��}!�V1� RQ��LIMIT_�a椀�M��CLmd}�R�IV	�a��EAR6��IO*PCC���2��B�Bg�CM@����R �GCLF�G!DYM(/�aR#5TWDG��| �s% �SS& �s>C P�a�!r1��wPQ_�!�(�!1��E�3�!3�+5�&�GR)A���?w��kP�W��ONT��EBUG)S&2*�p{@a�_E @ �p|�P�@�TERMB5�AK5ave�OR�IG0BK5sav��SM_�Pr�G0C~K5ved�TA�9�D�9UPB�E�3 -zAa�@.PY3>.@A$SEG�:f �ELEUUSE�@NFI,��2�1ޠ<p4�4B$UF6P��$�FQ4@��wAG0TQ�&�HSN;ST PATm�p�iBPTHJ�AߠE �p��2�P؀	E)�؁���1R�@�InaSH�FT_��1oA�H_SGHOR ܣ�6 �0�$�7�@Dq�'�OV�R#�na�@I�@�Uz�b �QAYLO=�z��I'"�oAj�!�j�ERV��:Qh��J ��OG @�B0����U>����R!P"�ASY1M.�"��1WJG�т�ES�A�YvR�U��T @���E)�ᥳEP�!�WP!�WOR @M|B��GRSMT��F�GR��3laP�A.@��p�q�uG ׸ ����TO�C�1�`P�@ �$OP��ဝpՓá �e�O��RE�`�RC�AO�pтpBe�`RmE u�h�A���e$PWR�IM�ekRR_�c4��qB� H2H���p_�ADDR��H_LENGqByqnq�q�uR��S�I H��S���q0Ӧu>Ӵu����u��SE�'�LrS<��J $J��`���_OFF��rP�RM� ^�aTTP_�H�wK (^pOBJ?"lip��$��LE`C�!�ȠL � \�׬�AB_~TS�bs�S{`��*�LVN�sKR��eHIT��[BG��LO�qt��fN�͂���`���`SS{ ��HW��A��M�p`INCP}U�"VISIO� ����+��t,��t,���� �IOLN��N�̠�C��$S�LQb��PUT_&�$�`{�P ��V���F_AS�"O��$L��I����A"��U�0�@Af��`q�<PHY���ÓZ�析UO��#P ` ������ڔ� �2�pP���`(�L��Y�,B�Z�UJ�Q�z�;NEWJOG-G���DISx�U�K�-�f�#R 
�WAV��ǢCTR�CǢFgLAG�"[�LG�d�S ���Y�3LG_SIZo����������FD)�I �4�E�*��D0�� �c$���𖶦���K��D0��� SCH_ ��߅p�2��N��F�T���E�"~���D����U
�
�{`L�n	�DAU/�EA�0-��dE�;�GH�b;�BOO��Uh3 Aɒ��IT��y��[0ŖREC��SC�R��ʑDIēS.@��RGO���˒� ���d�´���SU����W�Ĳ�Ľ�JGM�$�MNCH,�F�NKES0'�KM�PRGK�UFY�PYطFWDY�HL��STPY�VY�@Y؀�Y�RS��H1`uۺ�CT���R��� �$�U	�m���
R�ݠғ2`�G=��@POd����Ŧ�M�FOCU�d�RGEX��TU%IK�I{�����	�@�����I�M��@A��S�`���@������A�NA���2�VAI�Ll�CL!�UDCS_HI+4`�s_�Oe�
!h�S���|�9S����IGN4���F�J��T�be�_B�Uj � V !PT�$*��rv�ϤQ���a�!W !P�i�'���0�1?2�?3?��_� X � i�=a�5��L�Ņ�ID� tbP5R��bOh ��\A�ST�	�RF�Y� �@�  _W$E�C��y����^�� Y L�؟0��@�� �`qFtǀ�FwҬ�?_ Z �p�����b���>0C��[{ �p CLDP	�>�UTRQLI{��T8����FLG��� 1�O�D�����LqD���ORG�� ����hW>(�siT�r� 4\ �#0��Ք��Sy`T�70�#0' �$�!�#RCLMC�$B/T/�)Q��!r=1I�p_d] d��RQ73$DSTB�p�   6��-8�AX�R /8I<E�XCES�b�2Mp�1^�p2�T�2��0_�p"6_�A:&��;G?Y80K�d` \�GRO�U��t$MB �L�I9�CREQUI�RDB�aLO#KDESBUr� 1LYM���agbʑ`@�C�"F 1ND��`c`b��̨�CDC���IN'��C��Z`���H��N��a#�� �EP�ST�� c\rLOC�RITp��PAp�1 1OD�AQ��d X�O	N�cF�R�fV�	�X��b�U���uF�X0IGG�� e �y X�a��X4�XR�Q%��Y�	��X	��V�0ғDATA$`E�a��a��N��f t W$MDEaI:�)Sf��^d�![gH5P�@]exz��a_cANSW�aP^d�a��^eD�)AR�z�� Xpg �0C�U4�V�`�=URR2{�h D2�`A���A�! d$CA�LI&0��GS�w2NK�RINb�t<�'NTEg�(i�bCu���=RBqg�_N�qj@Pukr���$ht�2kuy7DIV�&DHi0jp:+�l $Vp�Cv�$�$Z0R�<!T 0R���b�em�H �$BEL�T˪ZACCEL���;�"�IRC�O�݁m��T����$PSi0�Lt� ڰW��Cp8��T�9�PATH���.���3]��Pl1_<�r���Ł�"S Cr��_M=G��$DD�9���$FW�`7`����.���DE�P�PABNe�ROTSPEEՂ@L� �JN�@��(0�t��$USE_p�P�&�ܦSY>��p�! ��QYN0A����OsFFua��MOU߁3NGJ�܀OL~�ٔINC�d2Q��-2x��� -2ENCSp�a2U��+4R�IN��I��B����"n�V�E��s^�23_UyPօp�LOWL��A[�` '���D>�@2@Ep]'��2C[p�W�MOS���4MO���0�'PERCH  ��OV����� �������$�8S+� � 2@������V�0^�O�L�P��7O�U��UP"�������TR�K��AYLOA �J��1����͵³3P� �RTI�1	�� MO�O�-2�28 �`4�wٳ��?�p�DUM2��S_BCKLSH_C�� P�ϐΦ����bn�"��y�Ñ���CLAL� V��!��� ��CH�K �SՐRTY@����C�
*!6a_�Nä_UM����C����SCL�W�LM?T_J1_L< 0-օa:�E4�U�G�pD�J�P�J�SPCd�0ȑZ���3�PC �3�!H_A@���C� csXT���CN_rN���.�S��%�V���:���ѹ�9�2��C' �SH�r �*�*!9�9� p��^����9���PA���_	P��_�"�Ŷ�0!ճ����JG�����~�OG��,�TORQU��ON��޹*�`B٢-�*�L�_W���_�sj��sj��sj�UIr�I��I�sFKP�]�J�!��c!�VC"�0'42��1��{08��82��JRK��+�� DBL_SMt���"M�@_DL�q�"GRVq�j�sj�sKH_��I���
�COS��LN - �����p�	�p�	 �����FZ� ٦�KMY�D�TH|�eTHET0��NK23�s��s� [CB�CB�sC&1�n2�����s��SqB�s��GTS�1W�C.�2Q�����$x�'3$DU�� �8A!r�2P&�19Qb8V$NE�4�PAI� ���"%�v$�p�A��%�'����LPH�5�"h��"S ��3�33�"+3(:2�pV�(V�(�p��,V�*V;V;V�";V0;V>;VL9H��(�&�2�-n�H;H�;H";H0;H>;H*L9O�,O�(O}I�.UO�*O;O;O";UO0;O>;O2F�"�Y�T�'SPBALANCE_T�@SLE�H_�S�PHq�hR�hR3PFULClX�R{W�R�3Uz1i
�UTOy_����T1T2�Y�2N���`��Tq@���Ps d���T��O�p!�L�INSE9G���REVf���Q�DIF��zy1jl_g�r1k��OBUa��t$yMI`���S?LCHWAR>���AB��u$ME�CH�Tˑ�a��AX˱Py��f�'�r�P�l 
�bI��:�ROB�CRW�-u��=)�pMSK_KP�t_n P �P_��AR��r_tn���18�c�a�_p`�y�_p�aI�N:a�MTCO�M_C���po � ݀g`4�$N'ORES��r��`�rop 8U�GRJ��eSD� ABג$XYZ_DA�!<F�r�DEBU:a�q����pq _P$��C;OD�� 1�����`��$BUF/INDXa�Hp"��MORRsr $�qU&���u��ӑy��W�!��bGi�s �� $SIMUL���8��>���F�OB�JEjP��ADJUySψAY_I���8�D���s�Ԑ_F-Iב=s�TZ�� c����`b�"�(�b`tp0G�D��FRIWÚd�Tg�RO%�A�Exb񊰓�OPWO> �Vpt0>�SYS�BU0[�$SOP���I�����U��b`PgRUN�rڕPArp�Dٖ�b��1�_OUbTΑ�a�t$�/IMAG��\pv �PDaIM��1�IN�[ �0�RGOVR!DY�˒���P�/�a�� L_�PB�}��¦�RB�� ��MLkᜪEDb��` �%N�@M��~���]��SLjPVpu x �$OVSLfS;DI��DEX���q �����o��Vb��N�A��'��,�'��D�M~�Ҥ_SsETK�Vpv @U�^��ep�RI��j�
Bq�_�}�����Hp�dà*� w Hx\q�`��ATUS<�$TRCx T�X�NѳBTMڷıI���P�4}Ѱ���Vpx D\pE���β�0�Ehbϱ�����ϱEXEհ����)�=��bf�ym�]p԰UP��L�$�`6�XNN����������� �P�G�uzWUB�ñ�e��ñ��JMP�WAI[�P���L�O7��pFA`��$�RCVFAIL_Cwq�p��R9��p�c���(�}�"�-�AR_{PL��DBTB��,��pBWD ��pUM*�"�IG�7��Q�c�TNLW�"�}�Ry�iӻ�E�����Hp���DEFSP` �{ L\p�`��_8��Ճ��UNI�����Ѐ�RD��Rb _L*A`Pͱ��P�pUq|-�#��q�O��XP:c�N�PKET�
���Pq�Uq} h~�ARSIZE5p���=��u�S̀OR~��FORMAT�P�g�COנq�<bEM2�d����UX��,���LIb�Uq~ � $�pP_SWiI�`��HqAXG�~b�AL_ o�J��A�rB���C�r�D��$EL����C_lі� �� � ���r��J�30 �r��TIA4�Z�5Z�6�rMOM���f��s���pB��ADf��s����PU�NR����s��������Rt�� A$PI�&E�kq E�p-~-�-��WC�0$��&��9q�gE��eSPEEDL@G�����Ծ ����)�9����)�8�	)���SAMWPx�p0�1��MOVD� H$_S`Y%nk%_��	1�t�2�t����c��v��8�H�PxIN ����������(�+(+GAMM�<Vu!�$GETHE�U�ٓD5�
�POLIBRv���I�$HIu�_L�ݰpB�&E�(A�.� �&LW�-�&�,�)	6�&�1��f�`j��� ?$PDCK���"ٓ_�����E� ��b7��a4��a9�� $I��R��`D�c�b~�Ե`L�E�qkq���81��0�pGq��`Vp�P/a?UR_SCR��A��r��S_SAVEc_D��8Ex�NO5�C��y�6�8@{$E�. {I��G	{I�@�J�KP �q��H� ���x" Mao���s���� d��6W2U�Cqy���:��M� �k�F� �aE��3�W<�@[�BjQWg@5r�U�R�R���Sc2jQM"��[C�L�W��M)ATr� ?� $PY����g$W`�fNG� O�`�b�b�b #�HЈ��a� ���c��%X�O���Z�e��ހRt� p䠰p�3+zO�O�O�O�O�a:5�_�r� |�E� 8@��>vs�>v��8@_��kwVvy�Eހu%\�(��"rB�\�P�"t�P���PM&�QU�5 � 8*�Q�COU�1 �QTH�#pHOL<�QHY�S��ESe�qUE��p.BZ�O��  bq�P���%��UNְ.�Q ��OE��p� P2�3��AÎ��ROG�����Q2�(�O}�2������IwNFO�q� #�he����RȾ�OI���� (�0SLEQ��с�рi�C�{�D$��L��`� OK0rj��!E� NU!���AUTTA�CO�PYqu�?��`@M"L�NI�M�X�Cᐛ�} Y�RGADJ�qe�i�X�Q��$�(���`��W��P���0��������EX8�Y%C0b�ѪObp�q����$�_NA9�!�������`���� � Q���P�OR�A�B�SReV0�)a�Y�DI��T_��{��������������5��6��7���8y���S8BL���m�MC_F�p��BPL9A8An�ȰR�� 9��Ѽ��$iB���n�d� ,�0FL-`LL�C@YN�[�M��=C?��PWRc��zL��!�DELA���8Y5�AD�a� ��QSKIP�� �Q�4�OR`NT2�Q ��P_4�� ַ@lbYp�� ��������Ƞ��ՠ���������9�1��J2R� L�� 46*�EXs TQ%�� ��(Q����p�����p����RDCf� �`��X9�R�p������r��A$RGEA�R_� IOT�2F�LG��vi��M%PC���B�UM_����J�2TH2N'�� �1�����G8 TN00 �����Ml��`I�8��REF:r1�q� l�h���ENAB{�(cTPE�0�1���i�m� ��^QB#��:��"������2�ҙ������P����&�3�Қ7�@I�[�m���&�4��������������&�5�Ҝ1�C�U�g�y���&�6�ҝ������P����&�7�Ҟ+@=Oas�&�8��������&�SMSK�q�|���a��E?A��M�OTEF����`a@��(Q�IOQ5��Ic(P��POW�0L�� �pZ�����#p%�L��U�"$�DSB_SIGN��1)Q%���Cl��S�232��b�iDEVICEUS�|,R'RPARIT���D!OPBIT`Q�Y�OWCONTR`;�(Q��O'RCU� �MDSUXTASK�T3N�p[0�$TAT�U`PU#�0L�����p_,PC9�$�FREEFROMqSp��%�GET�0��UPD(�A�2�V"P� J��� }!)$USA^����6���ERIO��P@bpRY�5:"_�>@ �P}1�!�6WR	KI[D���6��a?FRIENDmQ�P�$UFw���0T�OOLFMY�t�$LENGTH_;VTl�FIR�`-C��RSEN ;IUFI�NR]��RGI<�1ӐAITI��4G�XӱCI�FG2�7G�1��Ѐ3�B�GPR� A�O_~ +0!�1REЀ�E3�e��TC���Q�AV �QG8��"J���u1 ~! ��J�8�%��%m���5�0G4�X �_0)�L|�T�3H@6��8���%r4E3GU�IW�P�W�R�TD�� ��T��а��Q�Tm�{$V 2���H�1���91�8�02�;2/k3�;3�:iva �9=i�aa�^S�jRS$V��SBV�EV'�(V�BK�����&c �p��F�"{�@�2q�kPS�E��$.r8RC��o$AŠFwCPR��Gv]U�cS'�Ą 7���D3I�� 0�@qV`��p�d`A���E0�@��=�
B5�S!� ��aRHg����R�6�N SAX�!$�A�0L(A����rTHIC�1pY���h�t1TFEI�|�q�uIF_CH�3��qI�G�a�pG1@bxf���m���S@��7_JF��PR�ֱ��S��Ԁ�d ӎ$SР�Z�GRsOU�̃TOT�t�̃DSP�JOG����#��_P��"O������j��&KEPF(�IR����@M�R&@�AP�Qn�E^�`�!�[�SYS6��"[�;PGu�BRK�B �.��pIq�p��M���΂�`AD�!̃9�OBSOC׆�NӕDUMMY14�p�@SV�PDE_O�P�#SFSPD_WOVR=���C�L��OR�CNm0b�F.����OV��CSFR��pU���Fn���!#��C��A�"LC1H����РOV�s0���W�@M��ĥ:�R�O�#ߑ�_�p��s @@�u@VER�pns0OFSu@CV? �2WD6���2�ߑj2,Y���TR�!����E_FDOY�MB�_CM�D�B�BAL�b>�f��attV"Q �240/p��N�Gg�z�AMx�Z�0���¿�_M~��"7����8�$CA�7�D�����HBK81��I�O�5���QPPA�=�"�M�5�͵�~��DVC_DBxC�~� �3"�Т�!��1��糖�3����pЈ��*��U�3��CAB��2VӆPѣIP���c�O��UX�S�UBCPU�r	�S �P P���90^SQ׹c���."��$HW_AC�Т��S��cA�A~�pl$UNIT��}l��ATTRI"����	�CYCL��N�ECA��J�FLT?R_2_FI_�G(��9&�1LP�?�>�o_SCT�CF_��cF_��6��FS8!����CHA�1�w�8���"v�RSD�4"�����q�_T��PcRO��>�� EMy�_ܠ��8d��a 1d��a��DIb0!�?RAILAC��9RM��LOÐ C��Q�*q��3q���PRJ��SQ�pU�Cr�zs 	�FUNC��@rRIN'PѸ0���u��!RA��B �����F�Ğ�WAR�~���BLQ����A0��������DA����	����LD)0��Q�1�q��*q1TI�2rQǁ�p$xPR�IA1�"AFB�P�!|ߠ�<`�R����MOI��A�DFa_&@��51��LM��{FA�@HRDY�4ORG6 H���A�0| �MULSE&@x"�Q��a �G��	�����$dm$�1$1 ��|�0���� xm��EG�̃�`ARހ��09�2o���z�AXE�ROB��W�A��_�œS�Y������S�W�RI�@s1��SCTR�� ��(�E�ч 	%1��AB�( �/&�a�ӰOT�0^�	$ߠARAY�sf"���S@	��FI��*�$LI�NK���!�a_�%#�%{q�"X�YZ82�*�q�#OFIF���"�"�(j 	B�j�4С��n�3FI��%7�q���j���_J���%��#N�QOP_>$H+5�3F�PTB\1�2C�Цi�DU�&62�TURN��2r�5t!}��p��|7FL�`��Ӑm�0�%+*7�	� W1�. K�M��&82�Q�2rQ�#�ORQ��G��-(�+p���z�� 3q�E"��TF�GOV�@-A��M*��y�4�E:�E@�FW �J��G���D��o�*� � ��A7�P��y��E��A�GZU:ZU�CG�E)R���	6�E���B�TAFQ��)4����0r'�AXУa2 .q�c�W�c�W�c�W �p�Z�0�Z�0�Z%@�Z K@�Z��Z
!�V� �Y � 
i� i� *i� :i � Ji� Zi� ji� zi��a�iDEBU{�$v�u��;q��"F7O�n�AB��6��C9V�z� 
fr�� ��ukњw�!�w�!�w �1�w�1�w%A�wKA�w���\0��"3LAB"2|EwЄ�҂�3� O EERV�EN� � $nq�_NAǁ!_�PO����` f�M��_MRA��� d�  T���ER1R����~ TYi��R�I�V"0�S��TO	Q�T)PL��T�Ѕ�L�G�CJ �� p�PTl X���_�V1�b�Q���#�2B�2+�����/@��p��5�$W��V���5VN�[�$�@�⠲ �S���Q�	EHELL_CFGN߳ 5%�B_7BAS��SRvp0�.K� �S��J�ϐ1a�%Α2�3��4�5�6�72�8�RO���̌ � NL:�3AB8n��АACKwv���)�o�u0iႩ_�PU2�COq��OU��P��ӕ������TP�_KA1R�0��REm�� qP����QUE٩���@���CSTOPI_ALzs��� ��TĠ�� SEM�[�w�k�Mw�y�TYf��SO`��DI����Є�=�װ_TM>K�MANRQζ� �E��$KEY?SWITCH���찱�HE��BEAiT���EpLE����&�U��Fd�����SO_HOM� On��REF�@PRi�P�R� ��C@�O0�p ECO���� _�IOCM�4M�k������'�O� DH�!ۧH�U��;�M7x��@�3FORCߣf�� 􂰓OMq � @Etxk�U#Po1B�O�o�3B�4x��NP�X_AS��� 0�ݐADD��(�$�SIZߡ$VA�R�TIPr�q�G�A(ҷ��
�˨�r�t�n�SV�XC<����FRIF�R��aS%�7�x���NFѲ�EАO� x�PS�IڂTEC*�%CSKGL=�T�"�0&��V�D��>�STMTd
�o�P\�BW�@�?�SHOWw��P��SV� K�� ���A00�0�Q�� K���O���_���i���U5��6��7��8��9��A����6������20��F��
 �� ��U ����� ����0��� �J@��:�1G�1�T�1a�1n�1{�1���2��2��2��2���2��2�2�2� �2-�2:�2G�2�T�2a�2n�2{�2���3��3��3��3���3��3�3�3� �3-�3:�3G�3�T�3a�3n�3{�3���454��4��4���4��4�4�4� �4-�4:�4G�4�T�4a�4n�4{�4���555��5��5���5��5�5�5� �5-�5:�5G�5�T�5a�5n�5{�5���656��6��6���6��6�6�6� �6-�6:�6G�6�T�6a�6n�6{�6���757��7��7���7��7�7�7� �7-�7:�7G�7�T�7a�7n�7{�7ڈ�	��VP$�UP}D��  �Px���x�YSLO��� � ��հ�����QTAS�sTƠ���ALU}U����C�U��WFdQID_YLѳ�UHI�ZI�?$FILE_Σ�Tf�$u�_VSA��� h��+`E_B�LCK(�8bg�AhD_CPUQi��Qi����Sod_R1�ɢR ;��
PW,�d�[ �aLA�S��8�c�a�dRUN5��a �d�a�d��5��a�d�a��d �T�pACC����X -$&qLEN~�3t��&p䫠��Iѱ
�LOWo_AXI(�F1&q
�T2mwM��ɢ���I����Q�yTOR.�&p�{DW��s�LACE���&p�����_MAuйv�u�w�qTCV�|��wTڱ�;�1�<ѷt��H_��s��J����M��"ӠJ����u���u2q2��������s6�pJKцVK~��4���3ՃJ0����JJ�JJ��AAAL�����4�5Xr;�N1B�N���	��tL�p_k��'�*!q��� `5`GROU�PY�Ӳ}B$�NFLIC�����REQUIREv�EBUV�"q�����p2���#pɖ!qx�޳�� \��APKPRՐC���p
!�;EN�CLOz�,��S_M ���A��u
�!q��� 䣠M�C�r;�Xr|�_MGц�C��,`��N��pBRK��NOL述����Rϰ_LI���է����JޠѤP ��p��p���p;��pDD��p6�K��8����"q���� �ҒMr:ql�Gqz�PATHv�������Rxh�������pCNR��CA��է���INF%rUC�pwQ�Cd�UM�Yop�����Q�E:p�Gp�����P�AYLOAͧJ2=LHPR_ANqQÁL�`[�W�K�g���R_F2LSHR���LO\�䱕���>�ACRL_��ⵐ��޷C�XrH�P"��$H���FLEX�� qJ%u� :2Dv�p4�K�G`Yq�pPbt|F1K� �խ׃�������E����/�A� S�e�w�����y���ф����蘏����J�ÊT���X����υ �� څ��[����
�� � )��;�D�V�h�z�Y�}J��� � ��0�����QIPAT��ё6��EL4� �ؘ�J���ߐJE��C�TRޱ��TN��F��ɗHAND_V�Bp�ѹP`�� $&�F2��K��ШR�SWqX�j���O $$M��}�R���E��Uw�H��sA@�PH����Q���A���P��A��Aɫ���Tj`��D��DɫP��G�`1)ST��9!��9!N̨DY�`��� |�Y�鰋�KыǦ�@J�ч�s�U�ХP� �&�/�8�A�J�S�=��� ; �t�.Rx66N�/QASYM����Ґ����Խ��ٿ_SH�����筀�4��+�=�O�J�V��h�'CI����_�VI�dHN�u@V_UNI�ÉD���J҅�B�%�B�̦D�� �D�F�̓��������$*Uc���	Y���H�`��XQE�N� v�DIɠS�O�wT Y�YP��� ��I�1A��äQ �`Bc�S`�  p�a.a�� � MEB����R'R�1TkPPT�0) ���Qz�~�A��0�Xa	iT@�� $DUM�MY1��$PS�_��RF�ЈP$�Pf�aLA��YP��jb�S$GLB_T>mU�e�PpQ p8���Q� X	�ɗ�`�ST��ߐSB}R��M21_V��8$SV_ER��1OÐ�c�cCL�`�bEA5�O�RTPT O�P � D �`3OB���LO˰&u�q9c�`r�0�SYSqADR�TP�P�TCHb � �,&����W_NA����tz�9SR~���l = ��M�u`�ys�u~ �s��s������� ����0�)�T�"� 5�~���B����s�?�?��?D��XSCRE�)�p�ȐST�[�s}�P!��t�X�r _� Aq� T	��`ob��a`�l�P�Ҥ��g�c�O� �IS�c��TX�UE�T� �ñjp^`ySq�RSM_iq�mUUNEXCEPlV֑XPS_�a�����޳����޳R�CO�U�ҒS� 1�d�UE�tҘR�b9��PROGM� FLރ$CU�`POX?Q�д�I_�PH��� � 8џ�_�HEP�����PRY ?��`Ab_Ѹ?dGb��OUS�� �� @�`v$/BUTT�RV`��COLUM��U3��SERVx��PASNE� q��P@'GEU�<�F���q?)$HELPB�l2/ETER��)_�� m�Am���l���l�0`l�0l�0Q�INf���S@N0�� ǧ1�����ޠ �v)�LNkr� ��`rT�_B���$H�b TEX�*��ja^>�RELV��DIP�>�P�"�M�M3�?�,i�0ðN�jae����USRVIEWNq� <�`�PU�P�NFI� ��F�OCUP��PRI�a0m@`(Q��TR�IPzqm�UNP�T� f0��mU�WARNlU��SRWTOL�u���3�O�3ORN3�R�AU�6�TK�vw��VI͑�U� {$V�PATH���V�CACH�LO9G�נ�LIM�B����xv��HOSTN�r!�R��R<��OBOT�s��IM
�� gdS�P} 2�����a���a��VCPU?_AVAILeb��+EX��!W1N��=��>f1?e1?e1 �n�S��; $BACKLAS��u�n�\��p�  fPC��3�@$TOOLz�t$n�_JMPd�� ݽ��U$S�S�C6N�VSHI9F ��S�P`V�ȇtĐG�R+�P�OS�UR�W�PRADI��P�_cb���`|a�Qzr|�LU�A�$OUTPUTg_BMc�J�IM����2��=@zr��TILN��SCOL��C�� ��ҭ�Һ����� �����o�od5�?���Ȧ2Ƣ�0�T���vyDJU2��� _�WAITU���´n���%��NE>u��YBO� ��� $UPvtfaS�B�	TPE/�NEC��� �ؐ�`0�R6�(�Q��� ش�SBL�TM[��q���9p���.p�OP��MASf�_DO*�rdATZpD�J����Zp�DELAYng�JOذ��q �3����v0��vx��,d9pY_���9`7"�\��цrP? �N�ZABC�u� ���c"�ӛ�
�P��$$C��������!�PN�� � V�IRT���/� AB�Sf�u�1 �%�� < �!�/�/?? 0?B?T?f?x?�?�?�? �?�?�?�?OO,O>O PObOtO�O�O�O�O�O �O�O__(_:_L_^_ p_�_�_�_�_�_�_�_  oo$o6oHoZolo~o �o�o�o�o�o�o�o{|� ��AXLMT�vs��#  �t�IN&8qtPRE�O��+vupXuLA�RMRECOV ��)XrzujF ��%�!d�������7�I�[�m�~�,�� �/��uNG5� ��+	 =#��
ڏ�� PPLIMC5�?�%upՁ�Handl�ingTool �-� 
V7.7�0P/36 ���
]�_SW2�D�Fy0j�W� 43Y��J�9�K�7DA7�?����
&�X�e�	-�None���J����� �T7o�	�rP_��Viu�6s��UT�Oz"�,tTy.�HGAPON� %��!.��U��D 1�y� t�x�����y.��K�Q 1�{  THp������	��p�uq��"�"� �!��H�եw��HTTHKY��"ٯ���� u�����󿽿Ͽ��� ��)�;�M�_�qσ� ���Ϲ��������� %�7�I�[�m�ߑ��� �����������!�3� E�W�i�{������� ��������/�A�S� e�w������������� ��+=Oas ������� '9K]o�� ������/#/ 5/G/Y/k/}/�/�/�/ �/�/�/�/??1?C? U?g?y?�?�?�?�?�? �?�?	OO-O?OQOcO uO�O�O�O�O�O�O�Ƹ�TOĀ��DO?_CLEAND����{SNM  ɋ����_�_�_�_o��_DSPDRYR�_&��HI!��]@�_}o �o�o�o�o�o�o�o�1CU��MAX@ �bTQNQS�sqXbT�B�o�B���PLUG�Gb�cWo��PRC*4`B�P]klo^��rO�r=o��SEGF;�K�+�6��_�_�}�������ŏ�0�LAPZom�/��+�=� O�a�s���������͟�ߟ�6�TOTAL��v�y6�USENU
Z�g� HXL�NR���RG_STRIN�G 13�
��M,�S�
~��_ITEM1��  n󝬯��Я� ����*�<�N�`�r� ��������̿޿���I/O SI�GNAL��T�ryout Mo{de��InpB��Simulate�d��OutT��OVERRW` �= 100��I?n cyclHŕ��Prog Ab�or^Õ�>�St�atus��	Heartbeat���MH Faul<����Aler��� ��'�9�K�]�o߁��ߥ� ^S��^Q ��������,�>�P� b�t��������������(�:���WOR9���r���L����� ��������*< N`r�������PO���� ���9K]o�� ������/#/�5/G/Y/k/}/�/DEV� -�/�/�/ ??)?;?M?_?q?�? �?�?�?�?�?�?OO|%O7OPALT�� ^A��8O�O�O�O�O�O �O�O__(_:_L_^_�p_�_�_�_�_�_LOGRIxp��avO�_*o <oNo`oro�o�o�o�o �o�o�o&8J\n�_*�R�ݦqo ������(�:� L�^�p���������ʏ�܏� ���PREGbNK��$�r����� ����̟ޟ���&� 8�J�\�n���������~��$ARG_r��D ?	������� � 	$�	[�]���.���SBN_CONF�IG ��L��K�F�CII_S�AVE  ��k�b��TCELL�SETUP ���%  OME_�IO��%MO�V_H��¿ȿRE�P�|��UTOB�ACK��V�FRA:\8�� �8���'`��8�c�,�INI�a@8�^�,�MESSAGz�����|���ODE_D���}�C���O� ��,�P�AUS!��� ((O��J�\� F�|�jߠߎ��߲��� ������B�0�f�t��%�*TSK  �5ݒϕ�/�UPDT�����d����XS�CRDCFG 1v��� �������&�8�J�\�n� ��\�n���������� "��F��j|�����/e�2�G�ROUN����U�P_NAܰ��	�2��_ED��1�
��
 �%-BCKEDT-�0�}��p��ѲQ-2�p8�/�/�8���g2���E/��/��/~/��ED3n/&/�/J/�\.�/"?�/�/ED4 ?�/?�/\.[?�?5?G?ED5�?n?#O�?�\.�?jO�?�?ED6 ZOO�O6O\.�O_}O�OED7�O�Ok_�O�\.G_�_!_3_ED8�_�o�]-�_Vo�_�_ED9Fo�_�o�"o]-�o�oio{oCRoY_Vh�]1��{� LNO_D�ELGE_U�NUSE	LA�L_OUT �V��WD_AB�OR���~�5�IT_R_RTN�ǀH�ONONS)Ю������CAM_PAR�AM 1����
� 8
SONY� XC-56 2�34567890�Y �f�@����?�W�( С���8�h�х�ڎ��HR5ǃ��	���R570�B�Affފ������ڟ� ǟ�"���F�X�3�|����i���į!�CE__RIA_I����5��F��;�Я� ���GP 1]����s�����V�C󠸾�����CO�C ��(���ǀC8��@��H̺�CCX����Ch꺰p��x���� +C�����Ⱥ���+�=�G��ށ��HE>/pONFIG=�f��G_PRI 1�B�$r�����������(�~�CHKoPAUS�� 1���� ,wuj�|ߎ� �߲����������� 0�B�T�f�x����D�O���T���_MORGRP �2?� �\�� 	 �,��P�>� t�b���5�����eҒ.�?a�a�����K(���d�P�V��a�-`�/A�

s��������b&�i��ܦP�DB�����)
�mc:cpmidcbg��:�~�&��a���p�U�   �~�c
~�d3� ��d3�~��p.{C��e�/��/���{g�+/�n/�o�{f/s/i�u/�
D�EF �(K�)��b buf.t�xt�/�/��_MC�����z/2�3����ʇ�C�z  B�p�B��Z�B�X�B���~C� C�?��D3�u
q��Dv��D:�"�Df��ENN�EA7EV����=F�pgF=C��Fi�WG����Gp��G�/I�	ބ	6�����4���(D~*���/��ʄ3@9à1/  TB�D�V@2EI�5� F*� F��G$ˀF[� �GR�kNGl���G��G��&�H��G֓��H��߃]��  �>�33 �lށ�  N  ��@߂5Y�Ed��A���=L��<#�
 ��_�*~2RSMOFS���.^�9T1��D�E ��l 
� Q�;�P  x0_*_>TEST�")__��R���#o�^6C@A�KY���Qo2I��B�0��� �C�qeT�pFPROG %�(S�o�gI�qRu�����dKEY_TBL�  6��y� �	�
�� !�"#$%&'()�*+,-./01���:;<=>?@�ABC� GHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~�����������������������������������������������������������������������������q��͓���������������������������������耇���������������������9�Eъ`LCK�l��<�`�`STAT�c�_AUTO_DO���O�INDTO_ENB;���R�Q�Y�K�T2����STqO�~��TRL�`�LETE�ފ_�SCREEN �jkcsc� 	�UπMME�NU 1i  <�l�ol� K�u���FS����柽� ϟ���R�)�;�a� ��q���Я�����ݯ ��N�%�7���[�m� ������ɿ�ٿ�8� �!�n�E�W�}϶ύ� ��������"����1� j�A�Sߠ�w߉��߭� ��������T�+�=� ��a�s������� ����>��'�M���]� o��������������:#p)+�_M�ANUALӏ��DwBCOu�RIG��$�DBNUMLI�M�,1e
�P�XWORK 1k�_-<_N`�r�TB_� � m��Y0�_AWWAY��1G�@rb=�P�_AL� =���YҀ��`��_�  1!�[ , 

:&d2/(o/�&�Mt�IZP��@P�#ONTIM6��d��&��
�e#MOTNE�ND�o$RECO_RD 1'kU2)?�!�O�?1-?&k �k?}?�?�?88�?�? ??�?c?O*O<O�?�? rO�?�OO�O�O�O�O �O_�O8_�O\_n_�_ �__�_%_�_I_�_o "o4o�_Xo�_|o�_�o �o�o�oEo�oio�o BTfx�o�� /�����>�)� 7�t�� pu�����-� �͏ۏ�����N�`� Ϗ��o����)�;�� ����8���\�˟ݟ ����;�Q�گI���m���4�F�X��TO�LERENC�B��	"�L�Ͱ C�S_CFG (� +x'dMC:�\��L%04d.'CSVY� cֿx#[A ��CH�z _/x.�G��},���RC_OUT �)�- z/��SG�N *��"���#�17-J�UL-25 20�:52��2�7-MAY��14�:38�]� Z�t�����x.�����pa�m��P�JP��k�VE�RSION ���V2.0.�11~+EFLOG�IC 1+� 	d��ٓ���p�PROG_ENqB�2��ULS�'� �p�_WRS�TJN� ��"�E�MO_OPT_S�L ?	�]�
 	R575x#V?�74D�6E�7E�#50i�d�o�2E�d���j�"�TO  �.����k�V_� E�X�d�% �PA�TH A��A�\��M�_�~+ICTZ�F�, '�>`�eg��}��STBF_TTS��(�	��Eм`����� MAU��ߧ"MKSW��- )��},t���.�!��]l� R�v������4SBL_FAU�Ly�/��#GP�MSK�ߧ"TDI�A��0����`����!1234567890xS�l�P�����// %/7/I/[/m//�/�/��/�/�/L0PV ���/� 2?X?j?|?�?�?�?�? �?�?�?OO0OBOTO8fO8<x�UMP$�I�3 �ATR>㜢O�@PME���OY�_TEMP��ÈÓ3��4��DUN�I	�w�YN_BR�K 1��x�EMGDI_STA	����GUNC2_SC/R 27[��_ �_�_�_�&�_�_o o02or�nSUQ13y_+?�|o�o�o�olRTd47[�Q��o�o�� �_>Pbt��� ������(�:� L�^�p������� ?Ǐ ُ�0�,p��+�=� O�a�s���������͟ ߟ���'�9�K�]� o���������ɯ�� ���#�5�G�Y�k�}� ������ſ׿���� �1�C�U�g�yϋϝ� ׯ��������	��-� ?�Q�c�u߇ߙ߽߫� ��������)�;�M� _�q��ϧ������ ����%�7�I�[�m� ��������������� !3EW��{� ������ /ASew��� ����//+/=/ wa/s/�/�/�/�/�/ �/�/??'?9?K?]? o?�?�?�?�?�?�?�? �?OK/5OGOYOkO}O �O�O�O�O�O�O�O_ _1_C_U_g_y_�_�_��_�gETMODE� 15'Efa� t|�_GgR�ROR_PROG7 %�Z%���Ho�gTABLE  �[1O�o�o�o�Z�RRSEV_NU�M �R  ���Q�`a_AU�TO_ENB  qu�SZd_NO�a� 6�[�Q�b�  *�6p�6p�6p�6p�`+5pOastHIS�cXa�P�{_ALM 17.�[ ���6|6`+t���&�8��J�x_�bp  ��[4q�R���PTC�P_VER !��Z!6oZ�$EXTLOG_REQ�vs�y�SIZ�~܄TOL  Xa�Dz�r�=#�=
ނ_BWDo�%���fQ���_DI?� 8'Et�TXa< b[�STEPg�y�|�P��OP_DO�v�$v`FEATU�RE 9'EQ���QHand�lingTool� � DER �English� Diction�ary�7 (R�AA Vis�"� Master����
TE0�n�alog I/O���p1
0�u�to Softw�are Upda�teb� "/�k�m�atic Bac�kup
�d
!���groun�d EditB� � 25LC_ameraT�FX�� "Lo��ell�T��L, P��o�mm9�shۡ�h7600��cou����uct��p�pan=e� DIF����tyle sel�ectѡ- /�C�on��9�onit�or��Hd�tr~�ReliabT��ϣ(R-Diagnos��Q�	��H�Dual Ch�eck Safe�ty UIFc�E�nhanced �Rob Serv~��q �v	ԸUser Fr����T_i�xt.� DIO f�fiꫴ )�\�end�ܰErru�L�� ' prנ*�rO��� @���ENF�CTN Menurİv����.fd`��TP In?�fa]co�  
E�G��}p;�k Excذ�g�C��High�-SpeܰSki���  Par+�H����mmunicons��\ap���urf�?�X�t\�h8U���coknnZ�2Т !��Incr��str�)�8��M-6�K�AREL Cmd7. L��ua��}���B�Run-Ti.�Env�(<�@��I�<�+��s��S/�W�"H�Li�cense���� �ad���ogBoook(Sy>�m)	����"MACR�Os,��/OffKse\�f����H��!�Y�M1�Mec�hStop Pr�otZ�3� 5
��Mi4�Shif�\��B6S�Mi�xܰQ����H�Mo�de SwitcMhY�Mok���.�֥ ��Mt�Q�g�� ��5��ulti-�T������)�Pos�j�Regi>��� � ! �PA�t �Fun1��6iB9/��R�Num�Y��3�G�P/��� A�dju��	�/2H�S�)� o(�8�t�atu���AD n��RDMޱot��scove&� #�e�v�㱗��ues�t 867.��o��\���SNPX �b��Y���)�Libyr%�
�rt I��"�� "����.S�o�� ��s in VgCCM������ j�����㣀/Iހ� 710�TMILIBX�����g�Acc����C/=2�TPTX�� �Teln��Y@�����K�PCUn�exceptܰmotn�� �����~�\m725�����w�5���  h�640SP CSXC�i � j*��o RIN��We����50,��vrl�زmen" ��fiP-�a���P���Grid{�play F O/��? ̔�ELR;�|�20܁�ORDK�sc{iiw�load��41d�st�Pa9td��CycT�h�N��oriɰ:�7c oData� qu6�2�0�*�������7FRLamc�K��HMI De��(�����k�PC�φ�Password�7644��Sp������D#YELLOW� BO�	?1�Arc%�visu����#�ti�Op�^�! �2��aO�po�� t��ֶT1o�����3HT��xy�	��   $�t۠i�g��10Ơ 41�\+�JPN ARCPSU PR+��8b!OL0Sup�2fil� �!��E@-�;�croc�8�2��v���$ 12�jSS0e4�teex-� I�7�So�нtf�ssag�� �e��У�P��,��� {"Tc Virt���v�!����dpn��
�J3�SHA�Df0MOVE T��MOS O T�Ԡget_v�ar fails! l�>PU~1E����� Hold Bu�s %�h��VIS� UPDATE �IRTORCHM�A A�{�vYWEL[DTV S ]�DtS�: R741��o�uiPb}�y��BA�CKGROUND? EDIT "RC$�REPTCD C�AN CRASH� FRVR 62�z1�SCra��s �2-D��r ) �"��$FNO N�OT RE��RE�D �` m ��J�O� QUICK�aPOP FLEN� m41S�Loc<��gRTIMQ%�#�?FPLN: FG���pl m�r`�MD� DEVICE �ASSERT W?IT PCV;PB��AN#aACCESS M .pc��;Jo��Qui±��KbldmgUSB�$ ��t & re�mov�� Pg�S?MB NUL� ;a�|�FIX��C��AoCHIN,QOL�`MO OPT ՠ}a��PPOST0��WDU C�wQA�dd�`ad���0i�o�2��$P�`W�\0.$0`O�IN�&�P:fix C�PMO-046 _issueC�J/asO-�0�r130Т�- ��vRSET �VARIABLE�S-P{��R3D m~��view d���M��&�ea���b���of FD�5P�:N@x OS-1�y0`�h sc���t6��s t�lo��7 �WA�PZ�3 CN�T0 T�/"�I�mR�)�ca �Pu���POT:Whe�napewB�STYi E�{1t��ptKQdo GET_�p� �p��VMGR �LOl�REAd0C ~QW�~1�(�l�s�g�D�ECTpLpING IMPR�D�R(p+PB�PROG�RAM�ERIPE:STARTU� OAIN-;�ӠM/�ASCIIzPÂO�F Lq�DPTToB: N�pML$Gme P���`:x�;mo&�allW`!�.ӤTorc�A�U�dHC�iLpԸth�`n�@ ch��/GE�A�!�tou͐�R�Cal��k�Sig�n`� ND�ԗThresh123���`��09p : MS�G_P�+0er � �Q�Aܠzer�on��0 H85���RImA�n�2D���rc�0I��OM�Ea`�pONaP5� | נSREG:FF�-Д� ]�'���KAWNJI��n��J��9c�0asn d�!OA� immc �IN�ISITALIZ�ATI����~1we�m����dr+� L�B A�UWqmin;im�rec[�c!�R���m$�ro C-1>ѮS�ܰir�P�@ұJ�1pdETw��� 5`?�I�ow u���< se 1lc
��YbPM���p�Q��0�R`vR&�lu\�3ÏRe 0�4q�q1�#���m <a�ar�n��ঁBox �fo��*PRWRId�PW�S��v�09 �F�pup�de-�rel2 d�p� j���`━betwe���IND Q���igE snap|��us��spo T�ME��TPD#�D�O�p#aHANDL 1\k�`vR��Ȁ�D�ny�S�v�Yoperabil� ��T*�: H � l�\p��Vq�b�R�< p��a*�c&2O�`FA�,�.�-QV7. f�.v��GT�pib�s��� ɠtm�Line-Rem�ark �� RM�-�` W�#SPAT�H SA+PLOOS UIFc�+5f wfig�pGLA��D��Vrp������U�0�ther�V� T'rac���tW�\b�s7��d�t�� Mn�@  ���3:�ꕀdK�y��it �k8�d�PayR![�2]�ü1: g���s��dow�X�Q��0IS�q�qEM�CHK EXCE� C���MF +��Xah�� 35\!k��)���QBt� ��'b���[�c����e �`k�S�� B�UGr��cD$`PCETp���f�c4�~�0XPANSI���DIG��@OoPm�etTCCRG E�N��CEMENT4�A M̀K {�`�H GUNCHG9 �`� EXT�P�42�bQS�93 wP�8�x�ORYLEA=Kq  H5gyq��PLC WRDN� R �O /u�QS�PE=p��G*�V ���$�tn720\.3pGRI��A�r�T�PMC ETH���pSU7p�`  �j5/n�PENS�PN,��*P on=t�`BROW�`!sRMV ADDz 3CN qDC���P�T3 ALA2@ ����pSVGN E�ARLY�R��ŰH�57�GaJLA]YҀE (@M�P�PD�p*@H�S yI`P�OUCH8���V�F�q�com�H�x ��ERROR�� DE nJ��R=O�CURS8p�I��N4q�-1�58n7�RSR xP#aUp���Rqy�T�Fz�;�pk��Lt�� gՂ�B�SY RUNN��  a�`�BRK�CT�!RO�p3@ g\apSТ�AXxP����h8+ q��ISSUr} sPX�P�TSI�K1M1�0_�IPSAFE�TY Ck�ECK [��Á������<#8X�� �TWD2�@��@�INV��D ZOp�5X��t��DUALy� "MQ6�0�"rF#�E���dPdNDEX aF�t*UF�"�Pʀ�0sFRVO_117 A�PT6��KtqFALPTPW2477D6_�P�!n;HIG� CC�t�;SNPX� MM ��tq�d~�Vq�q�#�
"��DETEaC�Tq*@RRU��qA�P�5p�9 y�)�<9���7T��Pds� k�	��x�!Q���� t\4Ax�;A0�2 "Ke@" 8@HI�qXF8@4@�H�PRDC"�
@�aMB8@�IXF�b��� zOX@8@���a�G}E�B�Ccscr�J8@�Ndctrld.�A��NZE�A5��Q��!ĉ`�Df8@�`m�87�8�Q-;� ��� Krm`�
��PR̠78�@RI8@0q���Q (~\Mp��0t��!{B8@\tQ<OX�S�t0�3hB3nO�Vt9p�A�@LCF�L��{� �Rplcf��p�J8@�WTamai�E8@mubov2_miTA �O�S8@U`T[tT�AqP�r674xSSha?pe Gen��8@�j�I�[R�`�@8@T����%q (u8@��II�^�Q~C�a�[8@�;Ynrsg0�4� �3 4�CtMr68@�r�5hB5�zVnret-sp "r�Po�w{ng0bGCRE�pKa�ޠ�DAT�E��k�creat.��q�M�a�oksqg�tpad1P��(�tputZj�{�������܆28@����Q��f��sl�o��� �hexH�TB�8�ď��keyH�8@�pmZb�NR�u7A+�nrgc8@UQ�pp�bUZx�dp0aj921xSpl.Collأcq�\A��RNq�UA�3 (J�8@ip�_�W�A��_�Y��a7hB7��ͦtp[� "T�CLS9oKb��cl�skyh[��s�pkckZd���$�TQ����dA�rx�710a-� KAREL U�se Sp�FCTN9�a�7l�0s0a�� (���a��~C8@г�MI��c8hB8"�   �8@ �v	�v	 �  lmatea99�qM����E��mcclm5�CL�M;�� �j��E�et����aLM	�h�yas�p,���mc_mot�B�N��8@H����Q��su'��Q�ȕ������joi#�ߕ��A_log�Z����trc�B����ve��ϓ�v��QWX��6�f�inderxSCe?nter F1�lSw520��ha6rX� (<�r,�Q�Ձfi�Q �NH0�I�ۡ`���A8@uL��tq�a? "FNDRVϳ�~��etguid�UID�C8@������p���TA@�nuf;���P���ƞC�B��_z �Ӡo��qG������<l���fndrTY���2䁴tcp"�,qC�P MF�}38@5317��6s38�E ��gf6��(��K��Q`��-�X��A�tm6�P�İ��Q�`��	�͘��tm����b8@ej��TAiex��aP�Aa�ذ�cprm�A��l�_vars��
�� dwc7 TS��/�6���ma7AF�Grou�p| sk Exc�hangJ 8@�VM�ASK H5�0H�593 H0aH5�@� 6� 58�!9R�!8\�!4�!2���"(�/��;OMI� `@a0hB0�ՁU4U1#SK(x2�Q�0I�h��)�mq�bW�zR�DisplayImQ@vJ40�Q58aJ�!(P��;�� 0a��0��� �40;�qvl "DGQVL�D쌞�qvB�Xa`�uGHq�OsC��a�vrdq�O�xEscim�K40sJst]��uDdX@TRgOyB�B�v40)�wA~���E�E�asy Norm�al Util(�in�K�11 J�553m�0b2v�Q(lV40xU)������^��k986#8U����|�rP "NOR���dw d.a}oKksu �O�W���OY�W`�j0��6�H� menuu�yP6�M�`wRX�R5�77V�90 �RJ7989}�49b\:�`(�fity������e�<?��Vsmh`��8��C0�Sv�q��8���w�pn "MHMN<��ޣx �Ay`�o�3�u�`f�І�x�t��tRzQ��LV��vP�tm���|I�1{oPx �2|���I�y3I/B�odstǏ�ًmn����}enKsu_�L<���h!!���Rt��huseCrp��0Ҹ�ʐcM��_l�xP�oe��рpo�per����xdetbo/�l>�x����Ps$p�`���OPydspweb͓��z�'R��u�Rr101&S՟{t�`2�Z4�C30������`4�
�4�5��KQ�m[T��dUCalG40`�Q )p40}�����9;���DA�� v�	LATAumpd�\�bbk968��6�8c�fbl�4196�9y�9�|�D���b~d� "BBOX�|�M��sched��<��m�setuM:�����ff���40���n�41�ϒ�40q�co1l��|�1�xc�ؘ���li��X�0���j`��&�8�4 <�ro5�TP E�#��r�yK42r��;�(9T+Q �Rec'�� �1Iw�84�����Aok971��71�;����parecjo��QNS�[T���d�Xrail| naCgek�M ,QT2 *� (�ĜR%<�x�80!bh��p���4��4�yDgl�p�axrmr "X�RM�g�l�brf�{���n��kl��9turbsp��㧑�- �l015	�g�625C�Mh�+���@)89��	+��B6�� o�ҹ��x�7�q40�����pd "T�SPD�=��tsgl��l�:dQ����8Bct���K�vrE�aܮ�����?  �!����21�`( A�AVM �2�0 ��@fd TUP �him (J?545 l)�`8 �616 %�V�CAM ��C�LIO (�0�:�5&  (F\ M�SC �Rt"PBs�STYL�D!2�8 :2\ NRE �F2h SCH6p�DCSU tp�sh ORS�R �rD!04�S�EIOC& \f�xh 542 LE{X"� ESETn�X8!H ��sh8 7H ~�MASK��r�"7>��OCO*`	x�!03"6�!/40e0:66$ G639.6�[8LCH!6OPL�GR703
5MHC	R��0C� (! �0m6�A.f8!54
���00DSWb 58�8�180 �h!37 _88 (D�"02Cr24���27 q9�B25��2-6�05���9PRST ~bBFRDME�S�!zB�930 |_ NBA  6��� HLB 3 (�~!SM�@ Con>� SPVC �8!�20z��TCP �aram\T�MIL A��@PA}CETPTX �@�p TELN 9�6��29�%UEC�K��r UFRM� et�P!OR �ORP IPL%CS�XC�0j�1CVV�F l FQHTTP stA")�I#�� CGHP8Z�IGUI�0�hPPGS Tool� H8�@djZ��!@L�h!63�%�@32Q�\�31 B�h!96^�%R651�Rs�!53 TFAD�R�41�8"1 ��o�o�"9��4177�5�"/@�P�VCTO`�@�U�!sh!80�%�PRXY�R�!77�0 �b8 885 �ol3P� L� аdai� �`ڳh LCP<{Q� TSS �b�2�6:����@CPE :�HT@VRC~��tQNL ��@00�2 %��b	0dis� �`7 <��a\0�T��`1 �`en�b4� 652�`)FU0A2Q0Πo`p�Ptu�&r4 $r5N��R;U0p@nse�QJp?1 APFI[ Jp�3�g34�g40 �alxrE1t44�w46� ts UA0  7v�0O��r5�e��p7 p "sw&�a61:��r4��r5 QpwGr`�$�pQ8R�"sP`tQ�b��36w77�w8`�v8	3���r8�&:��pOq�8�8 "rkey�8�9F��a90�9�1 p�#@��� �D0�95�g97*pur�A1@d���P|P�q)1�0QplSq1p#4h��]a!s1@sl�B��8�Ӽ�\1�d1�`"��v�@{�14p�ae��5 h2��`�)6ޣ��7�f1p@��@d�YpCqd�ـd�1�`!uq��� Cu1< Oq4� ��7ReU1$ �u�1�Pϱ� ��@- �WQ158 as7e C��9 B��60 82ń�p�~��4 (Wai���`吢!��7E��86�EU1P`ro9�<�	1��<�2��<�	0����T��l�5J�l���cC���9%�MCR���P�2�`�Q2N@967�Q��8��
��9Z�2TPB���P�2P7U5@�o�İ�
�5�`U���3 �w���?A�E�1��c�qAwl��A�1��512 f��1�u5Р���a5p$��!56�+a��Q5h��҆��1 @��pp�b^[�538 xaB���|p�4�2�11/q5�p�4U5�P16 (߲�Pz��0��A8�P�����p�e5`��e5(�/�P`bbf�>�X��$Z�U�5d��\� X�7 	�  ��8 k_;kv��79 s�782 &�H5��E6���p����h���ñ����3J"�`��4 �3Ȥ59ѧ6�0t���8��6D0$�$�4 7��!���<��j670\tchk<�Ps��<�B<Ѓ90��7�<���<�\K�<�q�Ӻ�A�C<Р��q�<���<�t��sMg<�lc���FA<�H��<���<Я���<�hk��<Щ�B<� ��o�<���<��K�<�dflr��<Ш��� ��o�`���D�;�Z<�gEvam���� B<г�oќ���<а�|KЀ�creexl� ���P��<���|����j6<�s��prs.`���\���<�7��x����fsgn��P�b�t�at���<�L��1B !�svs�ch/  �Servwo S��ule>n�SVS��44�10u�_<��� (����/ched��,��~��A\�� �� B��@�B�qA����cj�+� � 5�1<����Ә�p�css "ACS<�&(��6@� �����c el����Q����tor�chms�<�- T��Ma`Ѵ���09� J5;598 �J681s�7� 8 ��b��<Чa����te,s�����8/�E�� m��wARC.�� 1q�a4�!=��C�tc�p�A�@t���f� F�����7#�2x�SE`�r���UtmSю0960'���RC������� p��96G= '��"H5W����L���\f�� �PATb����`!4U�#!Stmt�E ��� �pMA�!p��z�2?�in_<�X��r��X e/cW����pV����etdl��vߏ\oveto����܏��mmonitr�\��|#�0#st��?.6a��0PP���! Q�!�y`�`ame �Ar�ol�c�43�0a �p���01� �25�  ��<� v	��v	�A@�818\n; <s�I�B�2�pMPTP"��C�1mocol��,��C T�v�'!� �A���8P�53��y`Touc�hs�s�`��<��J5���Ѩ`mP����n[PQ�a,�E�a`��IP&
�Pth�A�<�KF#R�m;�Qet{th�THSR'��q-�Rt��o "P�GIO�#!$s�ISwka�"WK��!�MHqH54��5w5n/�Sm/��@ !7�*�da��8`!w�/Ac��tsnf T k�/�#gb�a��u`�
�^m�`u��Zӭ���Qp�є�#���Ka<��M��t5QtZ �a<��dFS5GK����G�1or��dW��64��tPx���P ����x,��?$���P�<�Z4e7�g "S�VGN.ox�copy "CO;�Wj$��O�A�9� "FSG@�ѧ�%7��_��f� �wQSWF*!"(�sgatuɀ���_
v��tp_TPDo��9�79�#dߎ?8���h�GAT���|!#��  �� �f�` ��"/� �w�Z� �b?6?� ����� ����E ���M� �ch�rT� �K6K� �sm�s� �o6�ѐ�gtdmen?3 �?��� �>��mkpdtd2 �0��, ���pdQ�X�� ����� ���mvbkup. �[�C�С���mkuno��p9rp���mkl �4��s �niU��� ��ldvrw���glg�4�� ��棑��7aut7�.pб����� �ַ������su 3� �Ǜ� �Ƿ� �2��\ �6�b2X� ���&�� �����A4��  ��B   946" ��fB� ��t\paic\p4k947 ���F#����� �ictas����pa`���cc�:�<��o�����geIn�� � ��F�lnpr � ����stf@��1��wbO�c��Ջ�8`��߄�vri�ߢ� а�-T� ���p��flow� OPAc���ow���R50�qtS �#T� (A���4�#���pѣV�c�u3�QF� ��SI�ac����46����s&��pa��!!���� ���55�b �o)��p���0娿
�afcal3�P� ��f��(}���`�f��m	߳� p�d�m�/���a/���$C`ѷ�� �! t�rack\P� 0�i�ne/Rail cTr�]TJ�69W�T  (L��8(`� �T.�`�%��D��P0�i (��8�48��_ɛ�⇒4����� �3�b3���3alV@ �NTf���%��Iin]0m���aen�������&?5�c@Itst3@��$����`� ,R9�%���0氱%���popener�s-OW dDev��F�M�6W���|A0�Pc"�l!esv� � ,��R��V$�Q���U<�LV$ �k9j �6���# �����%paop/!OPNU�V ��2celL��8�g_��/�6��ts�cG��$��V!�3� 5vrop�ߡ�7`�n(`�V"2D�a� V'O$:S9��� PumpE��jQ�@�"  ��!
��@бMSC#� @��)P��AC�`���� � v���� \mhplug�@!g�"7P��uK")���io7�CJ0��E讏LIO q1g 7�A93շ�5 q9� t����4rb ST��R��CPJ989�P�LSE�' �e eC3Q(P �/Ov�@���o�P� ? I1�R���55��f�I1�`�tcmio��McIO�����Utco1�"CL01V �c,BK`io��uM?���Sl�I0�ߢ�Eg �o���f �tI4\onfdtI���e%�p2�7�Inte�TB KCoMoo1E�R���(do554 (;r>Ex,��nR##�ipc�/>��qp5���
oQé�1�p�����7/o���ra�pd�CDV_��rP��8���qp2cnd��s
 �p��a�o�r`҄�S��"�c�a�c����2kIԿ?A�pcr!t���or0�qd#�� "���3p+���D��Џ��vr2k�0����AG�.+��cho�;�uC��(� �uV630�fwe P�m�����@���`��TX��� ��d�chp !"_��(	�3����p��8����\p3�v@����ш�9�3�1 �0����low�[�����chk���㳦As��s?Ө0�i�1h� ��2��i�w����s?1*�-	�:�O��vr������0�'����PFRAPWat?1rneE�P�sp�&� ac5� _A�rbo#�,�a��g���������Qs<�ICSP+ 9_����� ��F�A9P�H51IQ93 7���HX6hQ]PVR`S5���fPR6 iQWP�R� (P!am �S�u�"�A�I0�tpprg�0���`�h�@2atk932��!��E�^��asc �"8�C��S>i�atp�"�d�@1I�
g��dsblflt�JA�Qsable 'Fau�P{C!���EV0ex/!DSB (DC��t�$�p� �X 7� �� 5��Q��t3*�~���td9� "!%�(5��Csb9኏���\	��6#���@5�p$D@55�0-Adjust? PointO"tVJ�Rs�z�䐄��!�X�_�Yj��0\s�g��4��}7y�\a{da�"ADJ����j�Qetsha<�SHAP�sŭ'jpo�r4�t�!��@$ ��C|�	Tk!�bRPKAR/Qiagnostìy!O!vV66 J`(ew0�(�L��|�/�&krlde�  ��PP���hU b���r�3�Pp?q��DBG2C��� �X�o�1U�� ��WT�`�@ipJCM�aipper Opv`�1Se}78 (MH GF� ;":�&�##�� a�x�֕$��388C�����#�х9.�9C��g##PPk�Q��8�!�_"$�"�� =0%�P��A $��_�#%�0AQ�C~2 Mat?.HandlE��!�= &�pq MPLGET�0�1(�3�Tt& P�Sٰ'�B�1��B0� ���&p��H��PP �' p��@�C7PP	�TG��tD5�}m�q�Afh�nd "F_R  π����PP	 �  xT?Q���P(Pa��To�����?�pmpaO��JP^ ak925��2`H@O�JRpsQ`B2�u�nLHP�Tgse�GASo1�O�W�QT��0v !�R�Ptp~���JRdmon.�@��Vf�!ns�hYvr�Q J�g�Q�o�jY�HS~7�sl�f ��pen��PDnR(R&���ɐ823'��ٔq���g � ���� 1�� S�� ? �c\sltQ�!|Q E�P��a�rtPg��P��� �v��"SEDGp8�s0�qtdgY T����vP`ho �s`<`����qc�`g
�e` o�w�a@o"�'ile6�H�e�ȅ�nR�� �e! j�517�>Ճ��J@%��e�`��Q4��Q&�L�!F�J�=�ao�5�z/l17����_�œ��`C0C��  ��LANG j�ЁA��������g�ad���#�jp�.��4�Ē��ib���s�Ƒp�a���&���j5�39.f�,Ru~� Env
�������3H�z�J9�����h�Ф
Ҕ���2�2����� (KL�n-TiAmФ�⠤��p�3��TS����\kl�U�TIL"o���x�r "QMGl��!�8�����1 "��S��T3�\kcmn�o��SФT2���ut|�.�lreadc��}�exY�ܤ�r��\"��l��Фw�3��2C�*� -�C�D�E!�Ĥ� .��C� R C1V̴�Ҁ�\p�Р����p�tboxx��.�@�cycsL��:�RBTE�veriOPTNE���;ӕ�k�e�ߦ�a̸ߦ�hg�ߥ�DP=N��gp.v��r>�ptlit���0�4��te\cy�����tmnu�3`�r���5UPDT������8�駣��ite �� swto�,���oolB�F"�Y�`��Q��(q��gr3�@�䪒��"�䴁w������߳��s����� ��������lS���bx "O�� ����l����P���A�l\t�� ��������.	�Col�e!��R C��r��&r ��m;`��Chang��Lq�T1 �rcm 3�"��
� 6���"����sP7���"��222��2D2457�� CCFM�H���accda��Q�c ' ��KÕ0���K!����mo!���,$� ���!"
����/�/ ����	Y�,$��)�F,$sk����m rC%�tS1,$+��k1�%unc.,$oñ�1��sub������1��cce�5/!&��-/?-W/i&vs�}/�% #�#�/�.C��/� C%
�@? U �&+��F:q�t�
pDЃ D	  U�:7�~Dxmov.�P৅DPvc5Q�tfr�@PeC_UYgeob3dtg_y[tu���PH���PTUt�P�Sx�_r�^z�_�\var�_��\xy�_�[pclB`c�P���P�Ue�P?gripsuaosk�uti���ovfin�fpo}��o�j�b�P���Qud\�aX��P(c�\Rrp�Qnƅ�P�v�P)tm#qƆ�P�v�a+rog�a��\Q�?a+rpal?a{�{spa���P�u�Q�t�_�TZp�0�osipka�g3r�ovlclaAy(�:�t�pT�d�pu?a�c�A������ KtKa�P����qTf|�rdm��{rin#r���s� �2��b�|s�Pd�v�tv���v�h�0��ystn(* џ�yt'�1�p��aD�p�uϑ#�ul��@o�W6�2�siup1dl�]�o�vr�on��`1L�z�`\�r���gil3$|l4��ǉ#q54FyB�Տg{8�`���{wcmס����wxfer�UYt�lk2pp߿UYc�onv��sicnv�Qʯxag��H�Z�Glct`ao�=�p��׭nit0믁�3�x�����  ��� v	�v�	$��alϑpm�r&�B�eWa���f� %������I��߬�u�ͬ�KamT�f���c��w��roǁ#�5�����?� sm��y� a��y넑������`�����͐ϑ��p��m �Wa�1���A�6� S�e�X��ψ�\Q}��� ��������ĥw߉�� �߭���߮�#q0�� rs�ew���1�a��z긱n@�.�۲;�d�������  �> Ad	T$�?1 p! P��ve �e 	l�f@C�@�s/� � ?����8� ���<����reg.�C=~��o99 ~@�����$FE�AT_INDEX�  z ���e� IL�ECOMP :����1!�!z$#SETU�P2 ;1%~;"�  N f!�$#_AP2BCK� 1<1)  �)��/�/  %�/�/e4 �/�/>% �/$?�/H?�/U?~?? �?1?�?�?g?�?�? O 2O�?VO�?zO�OO�O ?O�OcO�O
_�O._�O R_d_�O�__�_�_M_ �_q_oo�_<o�_`o �_mo�o%o�oIo�o�o o�o8J�on�o ��3�W�{� "��F��j�|���� /�ď֏e������0� ��T��x������=� ҟa������,���P� b�񟆯�����K�� o�����:�ɯ^�� ����#���G�ܿ�}� ϡ�6�H�׿l����Ϡϝ���@)t Px/� 2� *.VR��߅�*�@߂�0F�j�T��PCrߛ�>��FR6:����V���z�T �!��K� ��q�S�G*.Fߢ��	��Đ���^����STM ��'���S����iPend�ant Pane	lS���HI���9���pU�������GIF�0;��������JPG��;��]o�R�
ARGNA�ME.DTy�">�\"���Rc�	PANEL1Y�%>��e�w��2�A/�//���/�3_/�/��/p/�/?�4�/I?��7?�/?�?TPEINS.XML�?�>:\�?t?�1Cu�stom Too�lbar�?Q�PASSWORDg?~w�FRS:\:O��? %Pass�word Config{OR��OSO�O �O��_�OB_T_�Ox_ _�_�_=_�_a_�_�_ �_,o�_Po�_Io�oo �o9o�o�ooo�o( :�o^�o�#� G�k���6�� Z�l�������ƏU� �y������D�ӏh� ��a���-�Q���� �����@�R��v�� ��)�;�Я_������ *���N�ݯr������ 7�̿޿m�ϑ�&ϵ� ǿ\�뿀��y϶�E� ��i���ߟ�4���X� j��ώ�߲�A�S��� w����B���f��� ���+���O������ ���>�����t���� '�����]�����( ��L��p��5 �Yk �$� Z�~��C� g�/�2/�V/� ��//�/?/�/�/u/ 
?�/.?@?�/d?�/�? �?)?�?M?�?q?�?O �?<O�?5OrOO�O%O �O�O[O�OO_&_�O J_�On_�O_�_3_�_ W_�_�_�_"o�_FoXo��_|oo�o�o�`�$�FILE_DGB�CK 1<����`��� ( �)
SU�MMARY.DG<�oblMD:�o*�n`Diag Summary+�8j
CONSLO�G qn�=q�Console �log�7kpMEMCHECK��2��qMem�ory Data|3�;g� {)�HADOW(������C�Shado�w Change�s���c-��)	FTP������=��qmment� TBD;�;g0<��)ETHERNET0�`n�q~����=qEthern�et �pfigu?ration��B`~%�DCSVRF/�p�'�@�C�%�� verify �allC��c1p=� �DIFF8���0�ůD�%Z�d�iffǯ{��q�1p������J� X��q�|�	�CHGAD�&�8�ͿD�ܯ�����2Ŀ����R�� `�yτ�GD �.�@���D�����FY3�ϳ���Z�� hρߌ�GD $�6�H���D�������UPDATE�S.$�
�ckFR�S:\"�c�>qU�pdates L�istc�`{PSRBWLD.CM���blN��e��pPS�_ROBOWEL \�6o+�=�loa��o�� ��&���J���n��� ��9��Jo���" ��X�|#� G�k�d�0� T���/�C/U/ �y//�/�/>/�/b/ �/�/�/-?�/Q?�/b? �??�?:?�?�?p?O �?)O;O�?_O�?�OO |O�OHO�OlO�O_�O 7_�O[_m_�O�_ _�_ �_V_�_z_o�_oEo �_io�_zo�o.o�oRo �o�o�o�oAS�o w�*��`� ��+��O��s��� ���8�͏ߏn���� '��� �]�쏁���� ��F�۟j������5� ğY�k��������B� ���x�����C�ү�g�v��$FILE�_N�PR]����Y�������MDONLY� 1<��U� 
 ��ۿ(���L� �5���Y��}Ϗ�� ��B�����x�ߜ�1� C���g��ϋ�ߘ��� P���t�	���?��� c�u���(����^� ������$�M���q�  �����6���Z��� ��%��I[���2����VIS�BCK����ų*�.VD�*� F�R:\V� �Vision V?D fileVd �������	/ ./�R/�v/�//�/ ;/�/_/q/?�/*?<? �/`?�/�??�?�?I? �?m?OO�?8O�?\O �?�?�O!O�O�O�O�O {O_�O!_F_�Oj_�O �_�_/_�_S_�_w_�_�o~�MR_GRPw 1=��Le�C4  B�`	� ��lo~li`���B��D���fnӺM�T� ��� ����e`i`a�o�khb �h�o�dcic.�N�pLn�eKك&M�7�GHD�E���|�i`@
��B���A�h�?
�7BX=��9�hl}A��[A�ZA���A�oA��T�pSl}F@ ��qhq�y�~g�fF�6�D�MqD��� BT��@���l}?pD���6���l����5��5���|��~e9�B��yA�bA�	ym�zsA-G*eA����z󏶈�����A�܏e�P����t�  @߬��?R�Z?AZ}@�r�{}�ޟɟ� �&��#�\�G���k�������zBH`� �����a;�Cީ���'�d
��Z��WZ����Q�HZ��@����@��33@����	\��[���ѿ�z�� 񿋯�*��N�9�r��]ϖρ�<�G�=��<�m]<��+=~�m<�c^��8eN�7��7ѷ�7�x7;��51���	ߤ��?߾dU2^`Yb`�b`��������F�`Үb` �b`��0����� C�^o�߂o�o�߸o� �o�� ]�(߁�l�� �����������#�� G�2�k�V�{������� ��������1  ��-�)��� ����0T? xc������ �/')�'/M/_/q/ 8��/�//�/�/�/�/ ?#?
?G?2?k?V?�? z?�?�?�?�?�?O�? 1OOUO@ORO�OvO�O �O�O�O��_��J��� �`_*�_N�_�O�_ �_�_�_oo'oMo8o qo\o�o�o�o�o�o�o �o�o7"[F jh�x�t�� !��E�0�B�{�f��� ��Ï���ҏ���� A�,�e�,/�������� �/�J����=�$� a�H�Z���������߯ ʯ���9�$�]�H� ��l�����ɿ��ƿ�� �#��O�OV� _z�D_ V_��z_�Ϟ_��� 
�C�.�g�Rߋ�vߛ� �߬�����	���-�� Q�<�N��r����� �����)��M�8� q�\������������� ����7"[Fk �|�|���� ֟3�WBg�t �����/�// /S/>/w/b/�/�/�/ �/�/�/�/??=?(? :?s?:�LϦ?p��?�� �� O��$O��T?]OHO ZO�O~O�O�O�O�O�O �O_5_ _Y_D_}_h_ �_�_�_�_�_�_�_o ��@o
�go*owo�o�o �o�o�o�o	�o- *cN�r��� ����)�;�M� ��������ˏݏď ��%��I�4�F�� j�����ǟ���֟�� !��E�0�i�T���x� ��ï�?�?��O��? OO�t�>O������ ѿ��ο��+��O� :�s�^σϩϔ��ϸ� ����� �9�$�6�o� 6o��Zo��R������� ���5� �Y�D�}�h� ������������� 
�C�U��y�����d� ����:�����+ Q8u`���� ���;&_ Jo������ //گ4/��x�j/4� �/X�n/|��/��/�/ !??E?0?B?{?f?�? �?�?�?�?�?�?OO AO,OeOPO�OtO�O�O ���O�O_�O+__O_ :___�_p_�_�_�_�_ �_�_o ooKo6ooo Zo�oZ��o�o�o�o�� xo
G2kR� �������� 1��.�g�R���v��� ��ӏ���	��-�� Q�/*/��N/��r/�/ ޟ�/��/)�D�M�8� q�\������������ گ���7�"�[�F�k� ��|�����ٿĿ���O �O�O��W�B�{�fϟ� ���Ϯ��������� A�,�e�P߉�t߆߿� ���ߪo��+�=� a��߅�p������ ����� �9�$�]�H� ��l������������� ��#G2W}h��p��$FNO �������
F0�� �  #�1 �D|�� RM_C�HKTYP  r� �q�� �� ���OM� _MI�N� m�����  X� SSB_CFG >� ~��Jl�Aj|�TP�_DEF_OW � m���IR�COM� ��$G�ENOVRD_D�O����TH�R d�d�_�ENB� �R�AVC_GRP s1?3� X� e/��/�/�/�/�/�/ �/�/? ?=?$?6?s? Z?�?~?�?�?�?�?�? O'OOKO2OoO�OhO��O�O�O�O�O�O�R�OU? E� �q������8�?#�O__K_m_�o_ꐖ  D3� ��_E�_q�@A��\Bȡ��R��>Y_6 WSMT<#FC-�U�foxo�o�HOST�C,1GY?ĭ�_ 	�h�k��o�f�oye CUgy�z1�������p	a�nonymous �5�G�Y�k�w��o�o �o������*� <��`�r�������ˏ 	�����&�8��� �����������ȯگ ���M��4�F�X�j� ����ݟ��Ŀֿ��� I�[�m�ρ�fϵ��� �Ϯ�����}����� ,�O�Pߟ�t߆ߘߪ� ����/�A�C�(�w� L�^�p����ϸ��� �������a�6�H�Z� l�~����������� 9� 2DV��z ������#��
 .@��������� ������//g </N/`/r/�/��� �/�/�/?Qcu� �/[?��?�?�?�?�? )/�?O"O4OFOi?�/��/�O�O�O�O9m�aE�NT 1H[ sP!^O_  `_?_._c_&_�_J_ �_n_�_�_�_o�_)o �_Mooqo4o�oXojo �o�o�o�o�o7�o m0�T�x� ����3��W�� {�>���b���Տ���� �����A��e�(�:����^�����㟦�QUICC0�̟ޟ?��1@��.�����2��l�~�߯!ROUTER௼�ί�/�!PCJOG�0��!192�.168.0.1�0	��GNAME �!�J!ROB�OT���NS_CF�G 1G�I ��Auto�-started^/4FTP:?� Q?SOBχ?f�xϊϜ� ���?�������+�� ��P�b�t߆ߘ�6� ����(�J� �1�C� U�g�6ߋ������� ��x�	��-�?�Q�c�  ?2?D?��������� )��M_q� ���:��� %t�����m���� ������!/3/ E/W/z{//�/�/�/ �/�/6HZ ?n/S? �w?�?�?�?�?�/�? �?OO<?=O�?aOsO �O�O�O�/
??.?0O _d?9_K_]_o_�_PO �_�_�_�_�O�_�_#o 5oGoYoko�O�O�O�O �_�o&_�o1C ogy����oT ��	��-�|o�o�o �o����o��Ϗ�� ��)�;�M�_�q���������˟ݟ�ÿT_ERR I������PDUSIZW  �^���$��>=�WRD ?�޵w��  guest+��}�������ůׯ��S�CD_GROUPw 2J� ��`�1��!��L_���  ��!��	 i-	�E����Q�E EATSWILIBk��+��ST 4��@��1���L�FRS:аTT�P_AUTH 1�K�<!iPendan�������!KARE�L:*���	�K�C�.�@��VI�SION SET���u���!�ϣ��� �����	��P�'�9����]�o޽�CTRL� L��؃�
���FFF9�E3��u���DE�FAULT���FANUC We�b Server��
��e�w���j�|���������WR_�CONFIG ]MY�X�����IDL_CPU�_PC���B��x�6��BH�MI�N'��;�GNR_�IO�K���"��N�PT_SIM_D�Ol�v�TPMO_DNTOLl� ��_PRTY��6��OLNK 1N�ذ�� 2DV|h��MASTEk��s�w�OñO_C3FG��	UO���>�CYCLE����_ASG 1O��ձ
 j+= Oas��������//r�NU�MJ� �J�� IP�CH�x��RTRY_CN�n� ���SCRN_UPDJ����$� �� ��P�A��/����$J23_DSP_EN~��p�� ?OBPROC�#��n�	JOG�1Q�� @��d8G�?� +S? /?)3�POSRE?y�K_ANJI_� Kl�H�3��#R�����5<�?�5CL_LF�;"�^/�0EYLOGG+IN� q��K1$���$LANGU�AGE X�6�e� vA�LG�"YS�߀�����x���i��@<𬄐'�0u8�����M�C:\RSCH\�00\��S@N_D?ISP T�t�pw�K�I��LOC��v-�DzU�=#�J��8@BOOK U 	L0��d���d�d��PXY�_�_�_�_�_� nmh%i��	�kU�Yr�UhozoLRG�_BUFF 1V��|o2s��o�R ���oq��o�o#, YPb����� �����(�U��D~/0DCS Xu] =���"lao�����ˏݏ�3n�IOw 1Y	 �/,����,�<�N�`�t� ��������̟ޟ�� �&�8�L�\�n����������ȯܯ�Ee�T/M  [d�(� :�L�^�p��������� ʿܿ� ��$�6�HπZ�l�~ϐϢύd�S�EV� ]�TYP�$���)߄m��1RSK�!O�c�"F�L 1Z�� � ���߯���������	�:�TP5@���>A]NGNAM�$�E���k�UPS PGI�|%�1�%x�_LO{AD0G %Z{%0_MOV�e����MAXUALRM;'�I(��~���D�#� V�#a��CQ[x�8��n��"�1060]\	 �F�	�� ��������������  D'9ze�� ������ R=va���� ����*//N/9/ r/�/g/�/�/�/�/�/ ?�/&??J?\???�? k?�?�?�?�?�?�?�? "O4OOXOCO|O_OqO �O�O�O�O�O_�O0_ _T_7_I_�_u_�_�_��_�_�_o�_,o��D�_LDXDISA�c���MEMO_{AP]�E ?��
 �5i�o�o��o�o�o�o�o��I�SC 1]�� �oTd��\no �������� �I�4�m��f���$� ��������!��E� ƏT�f�:�����ß�� ���z��ܟA�,�e� w�^������~���� �� �=���L�^�2� ��������߿�r� ��Կ9�$�]�o�(t_M?STR ^�͂ſSCD 1_xm� W���S�������=� (�:�s�^ߗ߂߻ߦ� ������� �9�$�]� H��l�������� ����#��G�2�W�}� h������������� ��
C.gR�v �����	�- Q<u`r�� ����//'/M/ 8/q/\/�/�/�/�/�/�s�MKCFG �`���/��LTA�RM_2a��2 �#\`Y>>G`METPUT`�"�����NDSP_CMNTs506��5�� b���>��"1�?�4�5POS�CF�7�>PRP�M�?�8PSTOL� 1c2}4@p<#�
aA�!aEqOG ]OO�O�O�O�O�O_ �O�OA_#_5_w_Y_k_��_�_�_�_�Q�1SI�NG_CHK  �+O$MODAQ�73d
?�7:eDE�V 	��	M�C:MlHSIZE�s0���eTASK� %��%$12�3456789 ��o�egTRIG �1e�� l��%��?   A$��ÜfYP�a,u���cEM_INF �1f>7 �`)AT&F�V0E0N�})��qE0V1&A3�&B1&D2&S0&C1S0=�})ATZ�� ��H�E��q9m��xA�u���X��������  ������v�)� ��я��П������� *��N�����7�I� [�̯ן���9�&�� �\����g�����i� ڿ������ï4��X� ��iώ�A���m����� ��߿�ѿB����� �ߜ�O������ߟߩ� ���>�%�b�t�'ߘ� K�]�o߁�����(� _�L���p�+�����������.ONITOR�0G ?ak   �	EXEC1T�#234Q5�`789�#��xx x*x6xBx NxZxfxrxU22�2�2�U2�2�2�2�U2�2�33��3aR_GRP?_SV 1g�y�a�(�Q?i=�?��vq��	@�M��
�y3<Hm�a_Di�n��!PL_NAME� !�5
 �!�Default� Persona�lity (from FD) �$�RR2� 1h)deX)dh�
!�1X d�/d/v/�/ �/�/�/�/�/�/?? *?<?N?`?r?�?�?�?�?�?�82S/�?O O 2ODOVOhOzO�O�Ob<�?�O�O�O�O_"_�4_F_X_j_|_�_LhRΐ 1m)9`\�b0 �_pb~�Q @D�  �Q?��S�Q?`�Qa�AI�Ez  xa@og;�	l�R?	 0`4bQ@4c.a�P�Jd�Jd��Ki�K��J���J���J�4�J~���jEa�o-a�@�x�o�l[`@�z�b�f�@�S��a��Q�o�c�=�N���
������T;f�
����m[`�*  �p�  �$p> p��$p��o?��?�������'���o�Bntr��Q�skse�}�l>�p�  �pu`�j  #p���vks�� 	'�� � �I�� �  ����}:�È6�ß�=���N��b@^�d��n�Q���{"�R�x���nN. ���  '���a�`@�a�@�t�@�p@p�n[`CpC�0�f0�+pB/pCz3}�P�@%��Ea  o�o$|m����gA%���. ����z�`�P���QD e���˟��(��m��� �t �O� ru �4 �R�<c��s� :	e�a��P�` �?�f�fd�!�����7� ��گ쬛af�F�>搠���iP�P�;�e�S�Ea4f�u��>LX��s�b<	��I<g�<#��
<2��<D��<��
vo��¯��S��S.���?f7ff?u�?&찗d�@T���?��`?Uȩ?X����Z���T:z�T B��Wa�з*dů�ρ� �ϥ��������&�8�0#�\�h�+�F. K� ��G߼�3���Wɯ�����G�@ G�� ��X�C�|�g�y�� ��������jZ���� ��Q����ߙ����� 3�������/A���t_�����������d���@+Fp�IP��t��%���[`B��0����<ze�xcb!@I�
��M`B@��@�`�9@y��?��h� �@��3�[N��N��N�E��<��/:/L �>���ڟ�A�p�C�F@�S�b/��X������@�t��%�h���`/qG���GknF&��FצpE,8{��/ F�ZG����F�nE�DE,ڏ�/�� ���G���F7��F��ED��.��C?.?g? R?d?�?�?�?�?�?�? 	O�?O?O*OcONO�O rO�O�O�O�O�O_�O )__M_8_q_\_�_�_ �_�_�_�_�_o�_7o "o4omoXo�o|o�o�o �o�o�o�o3W B{f����� ����A�,�Q�w� b����������Ώ� ��=�(�a�L���p������(r!3�ji̹�r���ꕢ�3�㱐ڟ�u�4 �����u�P�82�D�&�jb^�p��1w����� ����ʯ���ܯ� �Js�P^�PD�c�`� m���y�\������Ӱ�¿Կ�����.� G����}ϳϡ��� 홍�U�_�J���$�y.�@�v�d�z߈ߚ� x�4�������� ��D�.�2� �$[�G�[�^�B���B��CH� ^���� u����������p�h�M�_�q�������*���^�^�Y�rm�2��
 �� ��#5GYk} ������h*��� ��>�x}���$MSKCFM�AP  ��� ����m��N"ONREL  6�9_�"EXCFENBkq
7]�FNC��}JOGOVLI�Mkduyd"K�EYk�"R�UN��"S?FSPDTYU��<v_SIGNk}�T1MOT�z�"_CE_GRP� 1n��9\ ���/���/�/4��/? �/2?�/'?h??�?C? �?�?y?�?�?�?O�? @ORO	OvO-OoO�OcO �O�O�O_�O*_<_#_�`_-�"TCOM_�CFG 1o/����_�_�_
|Q_A�RC_�6��U?AP_CPL�_��NOCHECK {?/ 5� ;h9oKo]ooo�o�o�o �o�o�o�o�o#5�GTNO_WAI�T_LF'5y"NT��Qp/���q_7ERR�!2q/_�� R_���"��:�L�dT_M�O�sr�}, ���VP_��_�PARAuM�rs/���`���MW��� =e��345678901.�@�R�)�q���_� ����˟����ݛLW��3�E�؏i�cU�M_RSPACE�,�������$OD�RDSP�SI&�O�FFSET_CAsRToݨDIS��ݢPEN_FIL�E�I!�Q�v�POPTION_IO����PWORK 5t�'� T�|�/�^�F�U��Z����	 �m���C������RG_DSBL'  ��v����ޡRIENTTO�j��C���8=�#�?�UT_SIM_DJ�6	���VàLCT u��}\��Q��W�_P�EXE���RAT����� ���UP� ve������`�����*�8��$���2�#h)deX)�dh�O�X dY�ߑߣߵ����� �����!�3�E�W�i� {������������2n��)�;�M�_�q� ��������<��� ��+=Oas@���X��� O���1m(���(��.�g��"0 �дu�  @D7�  �?���?рH�D4  �EzZ3;�	�l	 0DӀS@SM� �i��i �H)!H�,�H8�H�m�G�	{Gǎ8��6�MV���� �C�)����)����Ճ�*�  �p  �z > �  ���/$"�,��B,�Btr�«�H�O¼�/���/��"�# �,0 �}� �  � �߽pj   ���&X�?MU	'�� � 12I�� �  ���-=���U?g;/�@}?�0~.ѱ�?�;Ѳ���H[N ��?A'M�D�> C%)�f)�" B& ��"O4B+�:�Q��@D1�oo�$�����JWAD0�J@�A: �1�E&?�O��O#__G_2]��� �t O�� ru �4� ��R�Uɳ�' :�%S�р�? �?�ff��@[�_�_V_{�o~��118р"o0j>�P�Q6YPрZo�WrAdS�%�>Lw0�#��<	�I<g��<5�<2��<D��<�ל���_��j�ѳMb�@?offf?�0?&p�:T@T�q?��`?Uȩ?X�-q�iyBq5Y a��gI�_� �����!��E� W�B�{���d�����Տ�LnpΏ/�ʈG�@ G��U�ȏy� d�������ӟ����� ��yB=� ��?p�� �/򏸯�߯R��� '�9��oN�`�����~�P����ۿƿ�B�� �D�e�ֿ;�ҿ_�J�?��h�oϨϓ�J���D4��b!�_@ ���� ߧ��Ŀ�����%�@I�)�M`�B@��@`��9@y��?��h	� �@�3��[N��N�N��E��<�/�Y�kЖ>��ڟ��A�p�C��F@�S���pX������@��t��%�h���߉!G��G�knF&�F׿�pE,8{�� �F�ZG����F�nE��DE,ڏ������G��F7���F��ED��Mf��b�M��q�� ����������(�� 8�^�I���m������� ��������$H3 lW�{���� ��2VAS �w������ /.//R/=/v/a/�/ �/�/�/�/�/�/?? <?'?`?K?p?�?�?�? �?�?�?O�?&OO#O \OGO�OkO�O�O�O�N=(]�3�ji�O�a���	U�E3Ա�x�O_<q4 ��%_<7_<q�P�Q_c_�ERjb}_�_1w?������]�Y��_�_o�_1ol��P�bPcn~���o�O@�o{_�o�oY�`��o �o,/;M#�f 0o�����Y�e@t�~�i#�1�C�yM� _�����������{bS� Ԏ��	�?�-�c�Mj�2���$�VG�Dz}�B����B��CH�}�9�֟��� ��0�B���wl�@~�������Ư�T�E��\��qQ��U
 ί�0�B� T�f�x���������ҿ����χ��� ���]{x}��$P�ARAM_MEN�U ?Յ��  �DEFPULSE��	WAITT�MOUTl�RC�V� SHE�LL_WRK.$�CUR_STYLvj���OPT��N��PTB����C��R_DECSNw� Te'�!�3�E�n�i�{� �߶߱������������F�A�USE_P�ROG %P�%�B��V�CCR���UeXÚ�_HOST7 !P�!����Tt`����������4���_TIME��� �T�  A�GDEBUG��P�V��GINP_FLM3SK]���TR����WPGA�� |�[����CH����TYPEM�Y�A�;�Q zu������ 
)RM_q �������/ */%/7/I/r/m//�/��/�/�/�/?��WO�RD ?	��	�RS��CPNeS�E��>2JO��ξBTE���TR?ACECTL�PՅ�Z� {`*/ +a`{`�>�q6DT QxՅ��0�0D��� #���0���2&��4'��Sc{a�0��B���5�0�2�0B�0@B�0��2��2�4U�4	�4�4�4�4�4�4 ��2U�4�4�4�4U�4�4�4�4Q�4��2�4�4���2!�4"�4�?�8 DOVOhOzO�O�O�O�O�O�O�O
Z%�9O.O @O2_D_V_h_z_�_�_ �_�_�_�_�_
oo.o @oRodovo�o�o�o�o �o�o_V!3E Wi{�����P���5�( �)� "�4�F�X�j�|�����0��ď֏��1u �*�<�N�`�r����� ����̯ޯ���&� 8�J�\�n��������� ȿڿ����"�4�F� X�j�|ώϠϲ����� ������0�B�T�f� xߊߜ߮��������� ��,�>�P�b�t�� ������������ (�:�L�^�p������� �������� $6 u�bt���� ���(:L ^p������ � //$/6/H/Z/l/ ~/�/�/�/�/�/�/�/ ? ?2?D?V?h?z?�? �?�?�?�?�?�?
OO .O@OROdOvO�O�O�O �O�O�O�O__*_<_ N_`_r_�_�_�_�_�_ �_�_oo&o8oJo\o no�oV�o�o�o�o�o �o"4FXj| �������� �0�B�T�f�x����� ����ҏ�����,� >�P�b�t��������� Ο�����(�:�L� ^�p���������ʯܯ � ��$�6�H�Z�l� ~�������ƿؿ��� � �2�D�V�h�zό��ϰ������$PG�TRACELEN�  ��  �_�������_UP y������������_CFG Mz�������<��� <�Z�l��<�$�DEFSPD� {/��a������IN'�TRLW |/���8L����IPE_CON�FI+�}����<�x�LI�D(�~/��GR�P 1���������@�
=�[����A?C�C�
�XC)��Bg��r�������dL�z������� 	 r�N��Ҩ掤� ´����B �����������A����> �6>7��D_������� ='?�=)����� ����	B-��Q��M���  Dz����
�� &L7p[�� ����/�6/!/�Z/��
V7.1�0beta1<��� B=q�"`�ff@��">�{���!=��͏!�A>ff�!@�f�f�"�\)�"D�_�?�  �!@�!L� �!Ap�#W��h/`??*?<?K;�w�����O/�?K/�?�? �?�?O�?O>O)ObO MO�OqO�O�O�O�O�O _�O(__L_7_p_[_ m_�_�_�_��_ o�_ $oo!oZoEo~oio�o �o�o�o�o�o�o �DQy{/�#F@  {yw}�y{ջy�-� �����/�Z?l?~? w���t�����я���� �����O�:�s�^� ��������ߟ�ܟ�  �9�$�]�H���l�~� ���_ۯ�����5�  �2�k�V���z����� ׿¿�����1�\n �j�|϶������ �	�4�F�X�j�c�� �ߙ߄߽ߨ������ ��)��&�_�J��n� �����������%� �I�4�m�X�����ί ����������!E 0B{f���� ��H�Zό�V h�ϴϊ�����  �2�D�V�O/�s/^/ �/�/�/�/�/�/�/?  ?9?$?6?o?Z?�?~? �?�?�?�?�?O�?5O  OYODO}O�O���O�O tO�O�O_�O1__U_ @_R_�_v_�_�_�_�_ �_"4FxBo|� ���o��o�o// 0/B/;�__J�n �������%� �I�4�F��j����� Ǐ���֏�!��E� 0�i��O^���N�ß՟ �������A�,�e� P�b����������o  o2oTo.�hozo�o�� ���o��Ϳ�o
گ '�֯K�6�o�Zϓ�~� ���ϴ��������5�  �Y�D�Vߏ�z߳ߞ� ���������1��U� ��y��:������� ��	���-��Q�<�u� `�r����������� T�f�x�n��� ��������� 7"[Fj�� �����!//E/ 0/i/T/f/�/�/�/�/ �/�/?�//?A?l�e? w?&?�?�?�?�?�?�? �?OO=O(OaOLO�O pO�O�O����*�O_�@RdZ_l_��$�PLID_KNO�W_M  ����A�TSoV ���P�[?�_�_ o�O&oo#o\o�B���SM_GRP 1���Z� dI`��oo$Cf�d_����D��T Pbj�oLk�f�o"~�U �o>n2T� ~�����7�4� ��p�D���R���ʏ ����������6�
�T�`�*������QMR�cń�mT�EGQK?  GR��(�#���[�� /�A�S����������� �$����W��+�=� O������������ �`��S�Ͻ�ST�a�1 1�����v�P0� @��� �E�ϲ��������� M�0�B�T�fߧߊߜ� ����������7��,�m��2�����A�<��z�3�������4���������A5)�;�M�_���6x���������7����������8(:L�ÿMAD  ����� ��PARNU/M  ��Ko����SCH�
 �
���S+UPD���xaq{��_C�MP_�`� <Pz '��U�ER_CHK����Z��ƪRS���_�Q_M�O� �%_��__RES_G����� ��v/{/�/�/�/ �/�/�/�/*??N?A?@r?e?w?J'��W,g/ �?L%��?�?�?N#(� �?OON#w�4OSOXO N#��sO�O�ON# �O �O�ON#d �O__N"�V 1��Uua�@�cX��Pp�P$@�cW،P��P@@�cV��P�"THR_INR���pbzA%d�VMASS�_� Z�WMN�_�SM�ON_QUEUEG ��e��`Ȩ`U�N�U�N�V�2`END4a6/Ni�EXE]oNeWBE�\`>o/cOPTIO�;g?+2`PROGR�AM %j%�1`O_�0bTASK�_I��nOCFG� �o�9pD�ATAɓ�B{@ev2w����� �z��+�=�O��s����������nzINFOɓ��}�!dr�� !�3�E�W�i�{����� ��ß՟�����/�@A�S�e�w�҇ބ��|� �98q�DIT� �Bׯj~WE�RFL~hwS~�RG�ADJ �ƪA�  ,�?E�8��Q~�IORITY�W����MPDSP(�a�j�U�WvT�;OG��_TG���R�j��TOE�P1��ƫ (!AF�PE5 ���!�tcp��%�!�ud�?�!icqm<�Q_��XY_<q��Ƭ�Oq)�� *������Op� �����������<�#� 5�r�Yߖ�}ߺ��߳�������&�*�POSRT�a�OpA%��_CARTR�EP~`Ʈ��SKS�TA�X!*SSAV�`�ƪ	2500H809u�T�T�䕣�ƫ������`X#�$�6�m�U�RGEU`B��A)W�FP�DO�V�2�W��q�?Q�WRUP�_DELAY ��Ưe�R_HOT��hwR%z����R_?NORMAL�n��<6SEMI:|y�QSKIP���X%�x 	 �������� X%-;%[mE �������!/ /E/W/i///y/�/�/ �/�/�/�/?�/?A? S?e?+?�?w?�?�?�? �?�?O�?+O=OOO1U�$RBTIF��>NaRCVTM�����m@DCR�����A;���BI�Y@�Y�?��ۧ�=�|����}`���uH�'_S<	��I<g�<#��
<2��<D?��<��
+__ {_�_)`���_�_�_�_ �_ oo$o6oHoZolo ~oi_�o�o�o�o�o�o �o DV�_z� ������
�� .�@�R�=v�a����� ������׏�*�m N�`�r���������̟ ޟ�����8�J�5� n�Y���}���ȯ��� ��A�"�4�F�X�j�|� ������Ŀֿ�ӯ� ��0�B�-�f�Qϊ�m� ����������,� >�P�b�t߆ߘߪ߼� ���������(�:�%� ^�A����ϸ����� �� ��$�6�H�Z�l� ~���{���������� �� 2Vh�� ������
 .@R=O�s� ����/�*/</ `/r/�/�/�/�/�/��/�/??&?28�AG�N_ATC 1���K AT�&FV0E02;�ATDP/6/�9/2/9p8A�TA2>,A�T%G1%B96}0k9+++�?�,�1_,�AIO�_TYPE  �EC/4?REFPOS1 1� K� x�O[H /O/�O�MNO`O�O �O�O_�OC_�Og__xd_�_+K2 1� KLON_�_o�_*o�_5A3 1��_�_�_� o�o�o�o@oS4 1�Woio{o�o3|W�oS5 1��o��oJ���jS6 1������]�H����S7 1��(�:�t��ݏ�>��S8 1������Ϗ	���r���)�SM�ASK 1� O � 
���ɗXNO��?���1.�8�1AMOTE  �.DN�_CFG �U����5�0BPL_RA�NGQ�K!Y�POW_ER �Q5 �a�SM_DRYP_RG %�%R����ȥTART �����UME_P�ROׯ�d�.D_E�XEC_ENB � �5]�GSPD�=����Y3��TDB̢���RMÿ��MT�_ѐT��S�D0O�BOT_NAME� �S�;9O�B_ORD_NU�M ?��A_H80�0I$��	��s	�\점��� ���e��	@�}�D|���D0PC_TIMoEOUT�� xD0oS232n�1�Q;� LTEA�CH PENDA1N��j�5��=Q��x0Mainte�nance Co#nsK"-��"+�t4?KCL/C�}��6��|� ?No Use�=[�8��F���NPO�ќ��5�_���C7H_L@��U����	J��MAVA#IL`���+��]�I��SPACE1 2�=L ����p��扢J@����8�?��� � ��V�w�N������� ��������4�&G 
l�}d	Q5U1��� ������`4&G�
l}d�#��2�������� 2A/b/%/w/�//�/�3����	/�/ -/O/^??B?�?�?�?�?�4�/�/??&? �?J?l?{O�O_O�O�O�O�O�5�?OO1O CO�OgO�O�_�_|_�_�_�_o�6_*_<_ N_`_o�_�_�o�o�o �o�o!�75oGo Yoko}o+�o�o��@��)��>��8R dv��H����ӏ%�F�-�[��Gw �� R�:;�
�� ���� ԟ���
��.�@�� ��c���p���8�¯=�dؠ��ϟ���!�3� E�W�i�_�q������ x��կ��'�9�K� ]�oρ�w��ϛ���Ͽ ѿ����5�G�Y�k� }ߏߡߗ��߻������� `S� @ ��8堯F�"�*ل�����߇��� ���,����V�h�2� <�N������������� .L4v�R@\n�����
f��7�_MODE � ��MS �"��&����Ïb�*	�&/�$CWORK_AD]���x�!R  ����t +/^ _?INTVAL]����hR_OPTI�ON�& h��$SCAN_TI�M\.�h�!R ��(�30(��L8�����!A��3��1�/X@>.?���S22�411d�8�1�1"3��@���?�?��?���IP���@���JO\OnOE@D���O�O�O �O�O�O__(_:_L_8O���4X_�_�_��8�1��;��o�� 1��pc]�t��Di�|1��  � lS2 ��15 17oIo[omo o�o�o�o�o�o�o�o !3EWi{� ���wc���	� �-�?�Q�c�u����� ����Ϗ����)� ;�M�_���`[���� ğ֟�����0�B� T�f�x���������ү������$�7�  0��� om������ ��ǿٿ����!�3� E�W�i�{ύϟϱ��� ����v���/�A�S� e�w߉ߛ߭߿����� ����+�=�O�a�s� �����ߖ����� � �$�6�H�Z�l�~��� ������������ `2DVP�\�  �A ������� %7I[m��������/ �/C(/N/`/r/ �/�/�/�/�/�/�/?�F;/?B?F��x1 ;?w=	�12345678�{��l�@�P�?�?�?�?�?O9/2ODOVOhOzO �O�O�O�O�O�O-/
_ _._@_R_d_v_�_�_ �_�_�_�O�_oo*o <oNo`oro�o�o�o�o �_�o�o&8J \n���o��� ���"�4�F�X�j� |������ď֏��� ��0�B�T�f����� ������ҟ����� ,�>�m�b�t������� ��ί����(��6yI�[�@�`����������Cz  B}p*   ����254F��$SCR�_GRP 1�(��e@(�l���0@} `1 [1�s	 )�3�C�<�t�vr�Y�8P�}�kϤ���[�95C����-�u��ȡ���L�R Mate 2�00iC �190��1Շ0LR2CA �3�=OÆ�D�
f؜1u�2�U7��`1��v��@�u���	t���������$�^0�2���_2T� gϡϊ��o�F�D�f?@��s�����￶ht �,Z�r�B�B˰�P�N�g�N�Aܰ�v�  @DЎ�N�@����  ?� ��J��H˰��y�N�F@ F�`������ A,Qwb�� �n�N�������B��_J �n�����/ �%//I/��E+:3��6?|?�5��
�/�/�#z��@=��"�/�pǢ� 3B�07Ƌ590@7���EL�_DEFAULT�  I����� ^1MIP�OWERFL  �V�v5]2�0WFD�Ok6 v5 �ER�VENT 1����O�t3C�L!�DUM_EIP�?�8�j!AF�_INEj0O�$!'FT�?=NOaO9!Q�O �PO�O�!RPC_MAIN�O�H��O�O�C'VIS�O�I��OE_o!TP8PPU<_��9d4_�_!
PM�ON_PROXY�_�6e�_�_XR�_�=�f�_)o!RDMO_SRV*o�9go�uo!RR8�o�4h,do�o!
�@M�_�<�i�o!RLSgYNC4y8�o>Y!ROS�?�|�4H�tO�8c� ����;��_�&� ��J���n������ ȏڏ7�I��m�4����X����7ICE_K�L ?%�; (�%SVCPRG�1�����!��3�*�/��4R�W��5�z���6�����7@ʯϯ�C��5�9��oG����o� �����D����l� �񑔯�񑼯7�� �_������4��� �]����������� '��տO����w�� %ϟ��M����u��� �������?�A��� ��ђ�؟ꐊ���ɱ ��������?�*�c� N��������������� ��);_J� n������ %I4mX�| �����/�3/ /W/i/T/�/x/�/�/ �/�/�/�/?/??S?�Ś_DEV ~�9�MC:[8�im4OUT�_Rf1~6i8REC� 1���f0�0} f0 	 f0]�2  
f0�4@�1���3OMK�1��4=A%O^OAA��
 ��Z�6 s;B�3AAqE=�=A���2WG�1f0)f0{�f0U�Of2B0��'���/Q0�O_��5��@��@r�H��;@�  x�0j}@U@��O f0)�f4�1af0�V_�2UX0��@�f0?�@��~_�__��2\J�0��0��0�@��[��_ f0�f0*�1=f0[f0�o�2UT0��@�f0*�@�u*oco�_�ÆLH��0�0��R ��  �RobmU��f0zf0�o�2�Q�*�@�f06�@z�oFvo~K�L=A�1(f0Etf0�f0�_c�f4�e�=�ZZ f0k�0��0Cf0f0q��"~N�LiI�1(�2�f2Pf0>jI�*�zDf0f0o.�g�V��φL"f0i�0Ubf0��0��0V��b�f0f0/f0|�~ 0��E0�
�@�f0$�@Y�^�p�
��ՆL*�A�0=�QpMɀ��b�ʈ��f0_^�f2C0��@��A0����&�C�2\�AM��Up#��A��p�<~��O���Ӧ�$2�k�ҟ��2\&f0}��0��0Wf0�Z��b�*f0f0R~�[���F%��@ݒq0"ޯ� *�a@��Z�H�~� l�������ؿ���� ��2� �V�D�zό�n� �Ϟ�����������.� �>�d�R߈�v߬ߚ� ���������*��:� `�N��f�x����� �����&�8��\�J� l�n������������� ��4"XFh� p������ 0B$fT�x�����5V 1�0�<��`!	O�2_ ��P��}�a?_TYPE�?�k2HELL_CFOG �z:f2/� HL�/<7RS ա�/�/�/"??F?1? j?U?�?y?�?�?�?�?��?O�?0OBOQK�
�p�!%QOO�O%���x�q�qQ��M�q�p�$�gBQ�d�O�O�&�HK 1��+ �OE_@_R_d_�_�_ �_�_�_�_�_�_oo *o<oeo`oro�oa&�#?OMM ��/�o��"FTOV_EN�M�t"!}*OW_R�EG_UI�o�"IMWAIT�b���G.${OUTv$&ywTIMu��`�VAL5's_UN�IT�c�v})MON�_ALIAS ?�e�i ( he !� ��$�6�%�� c�u�����D���Ϗ� ����)�;�M�_�q� �������˟ݟ��� �%�7��H�m���� ��N�ǯٯ������ 3�E�W�i�{�&����� ÿտ習���/�A� �e�wωϛϭ�X��� ��������=�O�a� s߅�0ߩ߻����ߊ� ���'�9�K���o�� ����b�������� #���G�Y�k�}���:� ����������1 CU y���� l��	-�Q cu�2���� ��/)/;/M/_/
/ �/�/�/�/�/v/�/? ?%?7?�/[?m??�? <?�?�?�?�?�?�?!O 3OEOWOiOO�O�O�O �O�O�O�O__/_�O @_e_w_�_�_F_�_�_ �_�_o�_+o=oOoao soo�o�o�o�o�o�o '9�o]o� ��P�������s�$SMON_�DEFPRO ����:�� *SY�STEM*  ��l�*�RECA�LL ?}:� �( �}Ecop�y md:cal�_dv_xy.t�p virt:\output\���over =>3�3030144:?694973�Џ�⏻p};z�frs�:orderfi�l.dat��tm�pback\=>�laptop-3�jv248ms:��48 ��G�Y��}2z�b:*.*��!�3�-�f�П���6x��:\�������P��B�T��7��a�@�+�2�ïկ�8z�~��v_z.ls~�@������D�V��Cz�z�����;�>�Ͽ� ����*���G�Y�l� ~�Ϣ�4�������� �� ���C�U�h�z�� ߰�6�����l�����ptcp.pc� ����D�V��5���_1ﱼ2�����h�z��2����F�X�����_��&�8������Az�ዿ�� +���Pbu���,� 3�������+� BT���ϔϯ�6 ��l�~ϙ�ϴE/ W/���Ϗ� �2/�/�/ hzߋ/�/���/G?Y? ����0?�?�?�? x�/./?OQOcO� O#O,/>O�O�Ot/? ?�/�OM___�/__ (?:_�_�_�?O�O&O �_Io[onO�Oo�O6o �o�o�O�O�_"_�oE Wj_|_2�� h?z?�?�?�A�S�e� x�����6�Ǐُ� ��"���E�W��_�_ o�2�ß՟hozo�� �o��A�S�e��o�� .��ѯ�v����� ��O�a�t������<� Ϳ߿����(���K��]����$SNPX�_ASG 1��������� P 0 '�%R[1]@g1.1fϰ�?���%���Ͽ� �����6� �@�l�Oߐ�s߅��� �������� ���V� 9�`��o������ �������@�#�5�v� Y������������� ��<`CU� y������& 	0\?�cu� ����/�/F/ )/P/|/_/�/�/�/�/ �/�/?�/0??%?f? I?p?�??�?�?�?�? �? O,OOPO3OEO�O iO�O�O�O�O�O�O_ �O _L_/_p_S_e_�_ �_�_�_�_ o�_�_6o o@oloOo�oso�o�o �o�o�o�o V 9`�o���� ����@�#�5�v� Y�������Џ��ŏ� ��<��`�C�U��� y���̟���ӟ�&� 	�0�\�?���c�u��� �����ϯ���F��)�P�|�_�x�PAR�AM ������ �	���P���p�OFT�_KB_CFG � ����״PIN_SIM  �ˁ̶�/�A�ϰx�R�VQSTP_DS�B�̲}Ϻ���S�R �	�� &� CAL_TC�ŵ�Ͻ�ԶTO�P_ON_ERR�  �����PT�N 	���A��RINGo_PRM�� ���VDT_GRP �1�����  	 з��b�t߆ߘߪ߼� �������+�(�:�L� ^�p��������� �� ��$�6�H�Z�l� ~���������������  2DV}z� ������
 C@Rdv��� ���	///*/</ N/`/r/�/�/�/�/�/ �/�/??&?8?J?\? n?�?�?�?�?�?�?�? �?O"O4O[OXOjO|O �O�O�O�O�O�O�O!_ _0_B_T_f_x_�_�_ �_�_�_�_�_oo,o >oPoboto�o�o�o�o �o�o�o(:L sp�������� ��9�6�׳VP�RG_COUNT������d�EN�B/�_�M��鴖�_�UPD 1�	�8  
M������ �-�(�:�L�u�p��� ������ʟܟ� �� $�M�H�Z�l������� ��ݯد���%� �2� D�m�h�z�������¿ Կ����
��E�@�R� dύψϚϬ������� ����*�<�e�`�r� �߭ߨߺ�������\�YSDEBUGn��Ӏ� �d��"�SP�_PASSn�B�?4�LOG �V΅�� ����
�  ��� �
�MC:\`��a�_MPCf�΅����ҁ���� ҁ��SA/V �i���� ���SV�T�EM_TIME �1�΋ (J�>�F�3�� ��T1S�VGUNSɀo�'������ASK_?OPTIONn�΅�������BCCF�G �΋O� H�2!`;A�I� r]o����� ��8J5nY �}�����/ �4//X/C/|/g/�/�/ ��,�/�/ ?? �/�/H?3?l?W?�?� �?��0�?�?�?O�? &OOJO8OZO\OnO�O �O�O�O�O�O_�O _ F_4_j_X_�_|_�_�_ �_�_�_o�X�  o2o Poboto�_�o�o�o�o �o�o�o:(^ L�p�����  ��$��H�6�X�~� l�����Ə���؏�� ���D�2�h�o���� ��ԟR�����.� �R�d�v�D������� ���Я����<�*� `�N���r�������޿ ̿��&��J�8�Z� \�nϤϒ���~����� �"�4߲�X�F�hߎ� |߲����ߤ������ �B�0�R�T�f��� �����������>� ,�b�P���t������� ������(��@R p������ �$6ZH~ l�������  //D/2/h/V/x/�/ �/�/�/�/�/
?�/? ?.?d?R?�?>�?�? �?�?�?r?OO(ONO <OrO�O�OdO�O�O�O �O_�O__&_\_J_ �_n_�_�_�_�_�_�_ �_"ooFo4ojoXozo |o�o�o�o�o�?  0BT�oxf�� �������>� ,�b�P�r�t������� ��Ώ��(��8�^� L���p�����ʟ��ڟ ܟ�$��H��o`�r� ������2�دƯ�����2��P��$TB�CSG_GRP �2����  �P� 
 ?�  {���w� ����տ��ѿ���/��A�T�[��b�d�0 �p�?P�	 wHBHA�L�͌�>@�B   C����0�ˀ��ϟ�D���ͣA���x���A��T8$�9��6ff��f�e@P�C�ώ�@�f����C��ߐ߮ߴ� ����%��%�D�W�"� 4���j�|�������?Y�����	�V3.00s�	�lr2c��	�*2�*�O�A� ��ѳ�33P�d��� 8x�J�y�  �������T�JCFG -��l� o���+��������=K
%�K q\������ ��7"[F j������� !//E/0/i/T/f/�/ �/�/�/�/�/s���? ?(?�/[?F?k?�?|? �?�?�?�?�?O!O3O �?WOBO{OfO�O�OP� <��O��O�O�O0__ T_B_x_f_�_�_�_�_ �_�_�_oo>o,oNo Pobo�o�o�o�o�o�o �o:(^L� �����h� �� $��H�6�l�Z�|��� ��Ə��֏؏� �� D�V�h�z�4����� ��ҟԟ��
�@�.� d�R���v�������� Я���*��:�<�N� ��r�����̿���޿  �&��>�P�b�ϒ� �ϢϤ϶�������� 4�F�X�j�(ߎ�|߲� ������������B� 0�f�T��x���� �������,��P�>� t�b������������� ��&(:p^ ����t���� �6$ZH~l� ������/2/  /V/D/z/�/�/�/j/ �/�/�/�/?.??R? @?v?d?�?�?�?�?�? �?�?OO<O*O`ONO pO�O�O�O�O�O�O_ �O__&_\_�t_�_ �_B_�_�_�_�_�_"o oFo4ojo|o�o�o^o �o�o�o�o�o0B �oxf���� �����>�,�b� P���t���������Ώ ��(��L�:�\��� p�����ʟ��� ��_ �*��_�l�Z���~� ����į�د� �2� ��h�V���z���¿ Կ濠�
�����.� d�Rψ�vϬϚ��Ͼ� �����*��N�<�r� `߂߄ߖ��ߺ����� ��8�&�H�n�\�� �>�����x������ 4�"�X�F�|�j����� ����������
 Tfx�D��� ���P> tb������ �//:/(/^/L/n/ p/�/�/�/�/�/ ?�/ $?6?��N?`?r??�? �?�?�?�?�?�? OO DOVOhOzO8O�O�O�O8�O�O�N  PS� V$_R�$�TBJOP_GR�P 2��E��  ?�hW<RCS�J\��@O0WP�R@T^�P � ��T�T� �Q[R	 ��BL  �UCр� D*W[Q�_�_?�fffe:l�B �P�ff@�`�33D   $a�U3o>g�_�_po�l��P�e9<�bbY��?٪``$o�o�UA��gD�`$��co�Quz9��P�Aa�P@a���C�Z`Ep�o]�A6ffpu`aD/�U�h�͔r��~ �a�RieAq�`�q��!@9q�|�d&`%����c333D�\P8o���?�`?L�pAp[QB�b�k�}� ���z�� >�ffԁL���T�f�� fo ��Nw@�*�8�f� ��r�,���П��ȟ�� '����F�`�J�X���,��SC�Vء��	V3.00�S�lr2c�T*���TQ�� �E���E�A �E��E��3�E�iNE�!h�E�فEۑ��E�I�E���E���E�r�F�F��FM(F�5�FBFaO�F�\F"f�,�z  E�@ �E�� E�� �E�  E������ E����� �EȆ�Ԏ�ᆰ��� F   F�� F$ Fj�` F�@ F��P F�` 9��IR9�o��D�L�_ ��V���LQ�8TESTPARS�XUP�9SHRk�ABLE� 1�J[4�SDV�+� �0�V�VȡV�WQV�	V�
�V�Vȥ�QV��V�V�뱅�RDI��TQ�϶���������f�On߀ۊߜ߮�H���ކ�Sl�RS 0� ������������� #�5�G�Y�k�}����� ��������/]k�o�� *	�%�7�I������+�=�O؆�NUM�  �ETQ��PP �밆�_?CFG �����Q@<PIMEBF_TTq��RS~�;GVER�<Q;�R 1�J[
 8I�RP� �@5  ����� �//&/8/J/\/n/ �/�/�/�/�/�/#?�/ ?Y?4?F?\?j?|?{�_�h@R
<PM�I_CHANG �R �3DBGLV�Q`IR;Q�0ET�HERAD ?*�E;@�S �?�?xTO6V�0ROUTe!JZ!�D�OwL?SNMASK0HRS>AA255.�E���O�O8TOOLOF/S_DIq��5I�ORQCTRL C�s[���n]8]_ �_�_�_�_�_�_�_o "o4oFo�
�_Tofo�o�g�PE_DETA�IH3ZPON_S�VOFF)_�cP_?MON �"P�2�iSTRTCH/K �J^mO�b�VTCOMPAT��h;C�d�`FPRO�G %JZ%C?AL_TCP=�n�%QPLAYr��j_�INST_M�@ 2�|�g�tUSe]�orLCK��{QUICKME�0)�oroSCREF�3Jtps��or�a�f��2w�_{���Zy�ISR_GRP �1�JY �� 6�����;�)�_�M��8���� Y�������͕��� ��/��S�A�w�e��� ����ѯ��������=�+�M�s�	12?345678�����f�X`�1�Ћ
 ��}ipnl/�۰gen.htm������0�B�X��Panel s/etupF�}<��`�Ϫϼ����� u� k��*�<�N�`�r��� ��ߺ��������� �ߝ�J�\�n���� �I�?������"�4� F���j���������� ����_�q�0BT fx����� ��>�bt�����3�~UA�LRM�pG ?J[
  �*/ !/R/E/v/i/�/�/�/ �/�/�/�/??<?��SEV  ��n6�ECFG ���m�6��A�1 �  Bȩt
  =?�s3E�?�?�?OO +O=OOOaOsO�O�Gz1ʂ��k SΟ�O�H7Isv?}{�`(% 0?"_p_I_4_m_X_ �_|_�_�_�_�_�_o0�_3o�L� �M�O�AoI_E�HIST� 1��i  �(p ��,/�SOFTPART�/GENLINK�?current�=editpage,�t,1}o�o�'{�(�o�eme;nu�b955�`�o�u��(:L148,2 _XYd��� ����}_r_AZ������2�'C�M~69n�o� ��$�86�ŏ׏,68n��`4�����3�M��}3�q��	��-���J�6��71n�MVn�������í�)a�a)o� ��%�7�I�ȓޯs� ��������Ϳ\��� �'�9�K�ڿoρϓ� �Ϸ���X�j����#� 5�G�Y���}ߏߡ߳� ����f�����1�C� U����ߋ������� ��Я	��-�?�Q�c� u�x������������ ��);M_q  ������� %7I[m� ������!/3/ E/W/i/{/�//�/�/ �/�/�/?��/?A?S? e?w?�?�?�/�?�?�? �?OO�?=OOOaOsO �O�O&O�O�O�O�O_ _'_�OK_]_o_�_�_ �_4_�_�_�_�_o#o �_GoYoko}o�o�o�o Bo�o�o�o1? �ogy�����o ��	��-�?��c� u���������L�^�� ��)�;�M�܏q��� ������˟Z���� %�7�I�؟������ ��ǯٯh����!�3��E�W�Bz�$UI_�PANEDATA 1�������  	��}  frh/�cgtp/wid�edev.stm�c���ҿ����)  ri��.�Ip��F� X�j�|ώϠ�ϲ��� �������0��T�;� xߊ�q߮ߕ���������Bv�� �   - ���@�E�W�i�{�� ������6������� /�A���e�w�^����� ����������+�O6s�l��  ��������� 1C�g���� ���L	///?/ &/c/u/\/�/�/�/�/ �/�/�/?�/;?M?� ��?�?�?�?�?�?0? Ot%O7OIO[OmOO �O�?�O�O�O�O�O_ �O3__W_i_P_�_t_ �_�_�_�_Z?l?o/o AoSoeowo�_�o�o O �o�o�o+�oO 6s�l���� ���'�9� �]�D� ���_o�oɏۏ��� �#�v�G��ok�}��� ����ş,������ �C�U�<�y�`����� ��ӯ����ޯ�-��� ��c�u���������� �T���)�;�M�_� q�ؿ��|ϹϠ����� �����7�I�0�m�T� �ߣߊ���:�L���� !�3�E�W��{�� � �����������r�/� �S�e�L���p����� ������ =$a����}�r�����)�*�� Vhz��� �����.//R/ 9/v/�/o/�/�/�/�/��/?�������$U�I_PANELI�NK 1����  � � ��}1234567890_? q?�?�?�?�?�4��]? �?�?OO1OCO�?gO�yO�O�O�O�OYIY0�:�M��[0  S�OFTPART/�GENA1?CON�FIG=SING�LE&PRIM=�mainedit �OI_[_m_YJ_$_�M=wintpe,1@_�_�_�_�]�_ $o6oHoZolooo�o �o�o�o�o�o�o
2 DVhz��� �����.�@�R� d�v��� �����Џ�����M 0, m 9P E=Por?S�5�co:�{�^��� ����͟ߟ��'� 9��]�o�R����O�O �����Z1�/�%�7� I�[�m�`C������� Ϳ߿񿀿�'�9�K� ]�o��L���э͙�S �����������#ߒS ;�M�_�q߃ߕߧ�6� ��������%��I� [�m����2����� �����!�3���W�i� {�������@������� /��Sew� ���.���|� #G*k}`� �����/�1/ C/֤�͡�ۯ}����/ �/�/�/�/?�2?D? V?h?z?�??�?�?�? �?�?
OO�ϝϯ�dO vO�O�O�O�OE�O�O __*_<_N_�Or_�_ �_�_�_�_[_�_oo &o8oJo�_no�o�o�o �o�o�oio�o"4 FX�o|���� �e���0�B�T� f����/������� ��ُ���>�P�3�t� ��i�����Ο��O/� s/(��/L�^�p����� �����?ܯ� ��$� 6�ůZ�l�~������� #O5OGO�� �2�D� V�h���Ϟϰ����� ��u�
��.�@�R�d� v�ߚ߬߾������� ���*�<�N�`�r�� ������������� &�8�J�\�n������ ����������m�"4 ßXjM�q�� ����BT 7x������A� �//,/>/P/C�t/ �/�/�/�/�/�/o/? ?(?:?L?^?Ϳ߿� �?�?�?�?�? OO�? 6OHOZOlO~O�OO�O �O�O�O�O_�O2_D_ V_h_z_�_�_-_�_�_ �_�_
oo�_@oRodo vo�o�o)o�o�o�o�o *�oN`r� ����m�� &�8��\�n�Q���u� ��ȏ������"����?�?�{��$UI�_POSTYPE�  �5�� 	k�{��_�QUICKMEN�  ��j�����R�ESTORE 1�ו5  ��/
�2�D�h�mc�������¯ԯ w���
��.�@��d� v�������W���˿ݿ O��*�<�N�`�τ� �ϨϺ����ρ��� &�8�J���W�i�{��� ���������ߡ�"�4� F�X�j������� ��ߋ����y�+�T� f�x�����?������� ����,>Pbt ������ (�L^p�� �I��� //��oSCREܐ?�u1sc-�Wu2M$3M$4M$U5M$6M$7M$8M!��USER/ 4/F"�T. O#ksW#�$4��$5�$6�$7�$8��!��NDO_CFoG ؜�  ,�� ��PDATE� �)�N�one V��SE�UFRAME  �
��&,1RTO?L_ABRT7?���N3ENBX?I8GR�P 1�!��Cz  A��3�1�@�?�?�?�?�?FO�"OG:ېUx81g;MSK  {5�Ag;MN41%a��B%���O��VISCAN�D_MAXyEI��c8�@FAIL_�IMGy@f���#��8�@IMREGN�UMyG
�KRSI�ZyC,���$,~SONTMOUW0�{D�%�VU�#گc�� �P�2�FR:\�O �� MC:\�XS\LOG�VB@4 !�O�_�Q�_�o
�z M�CV�_�SUD1&0fEX9k
�f�wV��2ۜ��p(��=7��͓o��j�o �o�o�o�o�o�o �2DVhz��KP/O64_?S�0��gn6�uQ0LI Q��z�x�qV� �|fy@�w�� =	�xwSZV�~����w�WAI��DSTAOT ܛ;�@�_ď֏�$����EP1�2DWP  ��P G/����q��AP-��B_JMPE�RR 1ݜ�
 � � 2345678901������� ʟ��ϟ��$��H��;�l�_�q����LT@M�LOW���P�@�P_�TI_X�('�@M�PHASE  �53��CSHI�FTUB1~k
 <���Ob��A�g� ��w���ֿ������ ���T�+�=ϊ�a�s� �ϗϩ��������>�@�'�t�K�!��#ޛ:	VSFT1�s�V�@M�� �5ԯ�4 �0��UAȯ  B8���Ќ"�0p�����Ҫ��e@F��ME*�{D�'��\�q��&%�!�M�$i�~k��9@�$~�TDINENDcXdHz�Ox@[O��aZ���S����yE����G����2�����������RELE��y?w�^_pVz�_ACTIV���H��0A ��K��B#&���RD�p��
1YBOX ��-�놫��2�D�190.0.� �83��25	4��2�p��&��ro�bot�ԟ  � pN g�pc� �{�v��x���$%ZABC�3�=,{�� �;-!/^/E/W/i/{/ �/�/�/�/�/?�/6?�?/?l?!ZAT�� ��